module _8inAND (clk, rst, Input_1, Input_2, Input_3, Input_4, Input_5, Input_6, Input_7, Input_8, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] Input_1;
  input  wire [0:0] Input_2;
  input  wire [0:0] Input_3;
  input  wire [0:0] Input_4;
  input  wire [0:0] Input_5;
  input  wire [0:0] Input_6;
  input  wire [0:0] Input_7;
  input  wire [0:0] Input_8;
  output  wire [0:0] Output;

  TC_And # (.UUID(64'd605037363922927401 ^ UUID), .BIT_WIDTH(64'd1)) And_0 (.in0(wire_11), .in1(wire_0), .out(wire_3));
  TC_And # (.UUID(64'd775080814455257473 ^ UUID), .BIT_WIDTH(64'd1)) And_1 (.in0(wire_5), .in1(wire_1), .out(wire_7));
  TC_And # (.UUID(64'd4575697617722991793 ^ UUID), .BIT_WIDTH(64'd1)) And_2 (.in0(wire_13), .in1(wire_6), .out(wire_12));
  TC_And # (.UUID(64'd2432098132025369908 ^ UUID), .BIT_WIDTH(64'd1)) And_3 (.in0(wire_9), .in1(wire_14), .out(wire_8));
  TC_And # (.UUID(64'd2530776218021452677 ^ UUID), .BIT_WIDTH(64'd1)) And_4 (.in0(wire_8), .in1(wire_12), .out(wire_4));
  TC_And # (.UUID(64'd2185451904912195012 ^ UUID), .BIT_WIDTH(64'd1)) And_5 (.in0(wire_7), .in1(wire_3), .out(wire_10));
  TC_And # (.UUID(64'd1870741422461363137 ^ UUID), .BIT_WIDTH(64'd1)) And_6 (.in0(wire_4), .in1(wire_10), .out(wire_2));
  TC_Constant # (.UUID(64'd4449029974404667643 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_7 (.out());
  TC_Constant # (.UUID(64'd1286176350726851474 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_8 (.out());
  TC_Constant # (.UUID(64'd357729215358331031 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_9 (.out());

  wire [0:0] wire_0;
  assign wire_0 = Input_8;
  wire [0:0] wire_1;
  assign wire_1 = Input_6;
  wire [0:0] wire_2;
  assign Output = wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  assign wire_5 = Input_5;
  wire [0:0] wire_6;
  assign wire_6 = Input_4;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  assign wire_9 = Input_1;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  assign wire_11 = Input_7;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  assign wire_13 = Input_3;
  wire [0:0] wire_14;
  assign wire_14 = Input_2;

endmodule
