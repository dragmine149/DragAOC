module Day2Part1z_Attempt2 (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_Constant # (.UUID(64'd1726993617052590723 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFFFFFFFFFFFFFFFF)) Constant64_0 (.out(wire_45));
  TC_FileLoader # (.UUID(64'd3987767967543158583 ^ UUID), .DEFAULT_FILE_NAME("day2_modified")) FileLoader_1 (.clk(clk), .rst(rst), .en(wire_71), .address(wire_4), .out(wire_0_0));
  TC_Constant # (.UUID(64'd337803116546834142 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_2 (.out(wire_71));
  TC_LessU # (.UUID(64'd2415299641673726094 ^ UUID), .BIT_WIDTH(64'd64)) LessU64_3 (.in0(wire_68), .in1(wire_4), .out(wire_1));
  TC_FileLoader # (.UUID(64'd4235385288069024156 ^ UUID), .DEFAULT_FILE_NAME("day2_test_1")) FileLoader_4 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_4), .out(wire_0_1));
  TC_Constant # (.UUID(64'd1484234401691717814 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_5 (.out());
  TC_DelayLine # (.UUID(64'd2141883989358176841 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_6 (.clk(clk), .rst(rst), .in(wire_47), .out(wire_64));
  TC_Add # (.UUID(64'd3665390526026043059 ^ UUID), .BIT_WIDTH(64'd64)) Add64_7 (.in0({{56{1'b0}}, wire_25 }), .in1(wire_4), .ci(1'd0), .out(wire_65), .co());
  TC_Not # (.UUID(64'd2915069602117248147 ^ UUID), .BIT_WIDTH(64'd1)) Not_8 (.in(wire_1), .out(wire_41));
  TC_And # (.UUID(64'd4444366698480428793 ^ UUID), .BIT_WIDTH(64'd1)) And_9 (.in0(wire_3), .in1(wire_1), .out(wire_30));
  TC_Or # (.UUID(64'd1455535717111312185 ^ UUID), .BIT_WIDTH(64'd1)) Or_10 (.in0(wire_67), .in1(wire_30), .out(wire_39));
  TC_Not # (.UUID(64'd4292279915901693506 ^ UUID), .BIT_WIDTH(64'd1)) Not_11 (.in(wire_3), .out(wire_67));
  TC_Switch # (.UUID(64'd259253643073170517 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_12 (.en(wire_41), .in(wire_21), .out(wire_8_1));
  TC_Counter # (.UUID(64'd4027361701724138616 ^ UUID), .BIT_WIDTH(64'd64), .count(64'd1)) Counter64_13 (.clk(clk), .rst(rst), .save(wire_57), .in(wire_12), .out(wire_12));
  TC_Ram # (.UUID(64'd3231836939472590219 ^ UUID), .WORD_WIDTH(64'd64), .WORD_COUNT(64'd1250)) Ram_14 (.clk(clk), .rst(rst), .load(wire_17), .save(wire_52), .address(wire_8[31:0]), .in0(wire_50), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_13), .out1(), .out2(), .out3());
  TC_Halt # (.UUID(64'd1646709671390234641 ^ UUID), .HALT_MESSAGE("Program finished!")) Halt_15 (.clk(clk), .rst(rst), .en(wire_63));
  TC_NoteSound # (.UUID(64'd2856162216424263791 ^ UUID)) NoteSound_16 (.clk(clk), .rst(rst), .command({{7{1'b0}}, wire_63 }), .note(wire_36), .pitch(8'd0));
  TC_Constant # (.UUID(64'd3448097267265053438 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h28)) Constant8_17 (.out(wire_36));
  TC_Not # (.UUID(64'd1023328388184503186 ^ UUID), .BIT_WIDTH(64'd1)) Not_18 (.in(wire_30), .out(wire_70));
  TC_DelayLine # (.UUID(64'd4092965687359902133 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_19 (.clk(clk), .rst(rst), .in(wire_65), .out(wire_48));
  TC_Mux # (.UUID(64'd316725708318265243 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_20 (.sel(wire_3), .in0(wire_45), .in1(wire_48), .out(wire_4));
  TC_Switch # (.UUID(64'd3903258603175327041 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_21 (.en(wire_7), .in(wire_13), .out(wire_24));
  TC_Switch # (.UUID(64'd1710097796709442780 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_22 (.en(wire_26), .in(wire_13), .out(wire_15));
  TC_Switch # (.UUID(64'd3052143593441878759 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_23 (.en(wire_38), .in(wire_14), .out(wire_8_0));
  TC_Constant # (.UUID(64'd3240501465042579115 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_24 (.out(wire_2));
  TC_Not # (.UUID(64'd1867582932362601439 ^ UUID), .BIT_WIDTH(64'd1)) Not_25 (.in(wire_57), .out(wire_28));
  TC_DelayLine # (.UUID(64'd2677504830674658084 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_26 (.clk(clk), .rst(rst), .in(wire_42), .out(wire_73));
  TC_Switch # (.UUID(64'd1725179244806057793 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_27 (.en(wire_35), .in(wire_24), .out(wire_42));
  TC_DelayLine # (.UUID(64'd1784992797701007900 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_28 (.clk(clk), .rst(rst), .in(wire_35), .out(wire_43));
  TC_DelayLine # (.UUID(64'd4350311000933170162 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_29 (.clk(clk), .rst(rst), .in(wire_26), .out(wire_9));
  TC_Switch # (.UUID(64'd4182440545682965520 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_30 (.en(wire_20), .in(wire_15), .out(wire_59));
  TC_DelayLine # (.UUID(64'd247377800554737393 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_31 (.clk(clk), .rst(rst), .in(wire_59), .out(wire_44));
  TC_DelayLine # (.UUID(64'd3700638478856170501 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_32 (.clk(clk), .rst(rst), .in(wire_20), .out(wire_56));
  TC_Switch # (.UUID(64'd3804153078929315197 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_33 (.en(wire_43), .in(wire_73), .out(wire_14_1));
  TC_Switch # (.UUID(64'd79719301686403854 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_34 (.en(wire_56), .in(wire_44), .out(wire_14_0));
  TC_Add # (.UUID(64'd1069550484725226130 ^ UUID), .BIT_WIDTH(64'd64)) Add64_35 (.in0(wire_10), .in1(wire_31), .ci(1'd0), .out(wire_27), .co());
  TC_Mul # (.UUID(64'd924182476717345043 ^ UUID), .BIT_WIDTH(64'd64)) Mul64_36 (.in0(wire_10), .in1(wire_31), .out0(wire_62), .out1());
  TC_Switch # (.UUID(64'd935510424511562668 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_37 (.en(wire_60), .in(wire_27), .out(wire_5_0));
  TC_Switch # (.UUID(64'd3389748284807452395 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_38 (.en(wire_22), .in(wire_62), .out(wire_5_1));
  TC_Halt # (.UUID(64'd3795677300099293191 ^ UUID), .HALT_MESSAGE("Opcode 99 Reached!")) Halt_39 (.clk(clk), .rst(rst), .en(wire_18));
  TC_Switch # (.UUID(64'd1224855048361981157 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_40 (.en(wire_40), .in(wire_5), .out(wire_50_1));
  TC_And # (.UUID(64'd4423175184107256786 ^ UUID), .BIT_WIDTH(64'd1)) And_41 (.in0(wire_19), .in1(wire_46), .out(wire_40));
  TC_Constant # (.UUID(64'd2201783711648500038 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_42 (.out(wire_46));
  TC_Not # (.UUID(64'd3940936562307563579 ^ UUID), .BIT_WIDTH(64'd1)) Not_43 (.in(wire_40), .out(wire_69));
  TC_DelayLine # (.UUID(64'd366563469061908473 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_44 (.clk(clk), .rst(rst), .in(wire_69), .out(wire_29));
  TC_Not # (.UUID(64'd23546066323564917 ^ UUID), .BIT_WIDTH(64'd1)) Not_45 (.in(wire_30), .out(wire_54));
  TC_Or3 # (.UUID(64'd1565632499214780517 ^ UUID), .BIT_WIDTH(64'd1)) Or3_46 (.in0(wire_38), .in1(wire_58), .in2(wire_70), .out(wire_57));
  TC_Not # (.UUID(64'd601742535760828746 ^ UUID), .BIT_WIDTH(64'd1)) Not_47 (.in(wire_51), .out(wire_23));
  TC_DelayLine # (.UUID(64'd1263282884327671549 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_48 (.clk(clk), .rst(rst), .in(wire_7), .out(wire_32));
  TC_Not # (.UUID(64'd4567426784455268513 ^ UUID), .BIT_WIDTH(64'd1)) Not_49 (.in(wire_32), .out(wire_61));
  TC_Not # (.UUID(64'd4522425577002129070 ^ UUID), .BIT_WIDTH(64'd1)) Not_50 (.in(wire_9), .out(wire_66));
  TC_Or # (.UUID(64'd571059853550174113 ^ UUID), .BIT_WIDTH(64'd1)) Or_51 (.in0(wire_18), .in1(wire_40), .out(wire_58));
  TC_FileLoader # (.UUID(64'd4032583951989155851 ^ UUID), .DEFAULT_FILE_NAME("day2_test_2")) FileLoader_52 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_4), .out(wire_0_2));
  TC_Constant # (.UUID(64'd1883781277529937826 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_53 (.out());
  TC_Constant # (.UUID(64'd4566527038733230091 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_54 (.out());
  TC_Constant # (.UUID(64'd3138890809031518109 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_55 (.out());
  TC_Constant # (.UUID(64'd2829021048917779791 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_56 (.out());
  TC_Constant # (.UUID(64'd1405985673201260239 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_57 (.out());
  TC_Constant # (.UUID(64'd3716163551666950261 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_58 (.out());
  TC_Constant # (.UUID(64'd4023943151529497828 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_59 (.out());
  TC_Constant # (.UUID(64'd2532988701438288488 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_60 (.out());
  TC_Constant # (.UUID(64'd4214058095318520776 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_61 (.out());
  TC_Constant # (.UUID(64'd958940107339709111 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_62 (.out());
  TC_Constant # (.UUID(64'd2113422115012713154 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_63 (.out());
  TC_Constant # (.UUID(64'd372203303927728035 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_64 (.out());
  TC_Constant # (.UUID(64'd4215445727210423365 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_65 (.out());
  TC_Constant # (.UUID(64'd4177145269316879433 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_66 (.out());
  TC_FileLoader # (.UUID(64'd3305349617174586722 ^ UUID), .DEFAULT_FILE_NAME("day2_test_3")) FileLoader_67 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_4), .out(wire_0_3));
  TC_FileLoader # (.UUID(64'd231382507668522051 ^ UUID), .DEFAULT_FILE_NAME("day2_test_4")) FileLoader_68 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_4), .out(wire_0_4));
  TC_FileLoader # (.UUID(64'd1231532553883646540 ^ UUID), .DEFAULT_FILE_NAME("day2_test_5")) FileLoader_69 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_4), .out(wire_0_5));
  QuickSave # (.UUID(64'd2695330121804011308 ^ UUID)) QuickSave_70 (.clk(clk), .rst(rst), .Value(wire_0), .\Number_(stored) (wire_68), .\Saved?_1 (wire_3), .\Saved?_2 ());
  BytesToNumbersz_3 # (.UUID(64'd1729469431074511873 ^ UUID)) BytesToNumbersz_3_71 (.clk(clk), .rst(rst), .Main_8b(wire_0), .Carry_In(wire_64), .Output(wire_47), .Offset(wire_25), .Value(wire_72));
  OnOrOff # (.UUID(64'd3163142382288365090 ^ UUID)) OnOrOff_72 (.clk(clk), .rst(rst), .Input(wire_41), .Output(wire_52_0));
  flippedzm64bzmswitch # (.UUID(64'd2031059029553199162 ^ UUID)) flippedzm64bzmswitch_73 (.clk(clk), .rst(rst), .Input_1(wire_12), .Input_2(wire_28), .Output(wire_8_2));
  OnOrOff # (.UUID(64'd150349705086353648 ^ UUID)) OnOrOff_74 (.clk(clk), .rst(rst), .Input(wire_28), .Output(wire_17_2));
  OnOrOff # (.UUID(64'd224193335304047014 ^ UUID)) OnOrOff_75 (.clk(clk), .rst(rst), .Input(wire_55), .Output(wire_17_0));
  mand # (.UUID(64'd3349436745291189726 ^ UUID)) mand_76 (.clk(clk), .rst(rst), .Input_1(wire_38), .Input_2(wire_2), .Output(wire_55));
  mand # (.UUID(64'd242248694494001734 ^ UUID)) mand_77 (.clk(clk), .rst(rst), .Input_1(wire_30), .Input_2(wire_29), .Output(wire_51));
  flippedzm64bzmswitch # (.UUID(64'd1881707450118815654 ^ UUID)) flippedzm64bzmswitch_78 (.clk(clk), .rst(rst), .Input_1(wire_24), .Input_2(wire_32), .Output(wire_53));
  OnOrOff # (.UUID(64'd4158355321388927517 ^ UUID)) OnOrOff_79 (.clk(clk), .rst(rst), .Input(wire_43), .Output(wire_38_0));
  flippedzm64bzmswitch # (.UUID(64'd558922318308219109 ^ UUID)) flippedzm64bzmswitch_80 (.clk(clk), .rst(rst), .Input_1(wire_15), .Input_2(wire_9), .Output(wire_11));
  OnOrOff # (.UUID(64'd3868852299644989347 ^ UUID)) OnOrOff_81 (.clk(clk), .rst(rst), .Input(wire_56), .Output(wire_38_1));
  Opcodez_zmz_1z_2z_99 # (.UUID(64'd1253066027045582023 ^ UUID)) Opcodez_zmz_1z_2z_99_82 (.clk(clk), .rst(rst), .Opcode(wire_33[7:0]), .Add(wire_60), .divide(wire_22), .halt(wire_18));
  OnOrOff # (.UUID(64'd779081389060044986 ^ UUID)) OnOrOff_83 (.clk(clk), .rst(rst), .Input(wire_40), .Output(wire_52_1));
  flippedzm64bzmswitch # (.UUID(64'd3330710435434371616 ^ UUID)) flippedzm64bzmswitch_84 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_40), .Output(wire_8_3));
  flippedzm64bzmswitch # (.UUID(64'd3395453474976780481 ^ UUID)) flippedzm64bzmswitch_85 (.clk(clk), .rst(rst), .Input_1(wire_72), .Input_2(wire_54), .Output(wire_50_0));
  CellWritter # (.UUID(64'd1760994904368207804 ^ UUID)) CellWritter_86 (.clk(clk), .rst(rst), .Clear(wire_23), .Write(wire_17), .Value_1(wire_13), .Value_2(wire_33), .Written(wire_34));
  CellWritter # (.UUID(64'd2225673571882546958 ^ UUID)) CellWritter_87 (.clk(clk), .rst(rst), .Clear(wire_23), .Write(wire_32), .Value_1(wire_53), .Value_2(wire_10), .Written(wire_16));
  CellWritter # (.UUID(64'd640733034693975124 ^ UUID)) CellWritter_88 (.clk(clk), .rst(rst), .Clear(wire_23), .Write(wire_9), .Value_1(wire_11), .Value_2(wire_31), .Written(wire_37));
  mand # (.UUID(64'd2253745888330672149 ^ UUID)) mand_89 (.clk(clk), .rst(rst), .Input_1(wire_7), .Input_2(wire_61), .Output(wire_35));
  mand # (.UUID(64'd4089700112481536660 ^ UUID)) mand_90 (.clk(clk), .rst(rst), .Input_1(wire_26), .Input_2(wire_66), .Output(wire_20));
  CellWritter # (.UUID(64'd3735606448599014512 ^ UUID)) CellWritter_91 (.clk(clk), .rst(rst), .Clear(wire_23), .Write(wire_49), .Value_1(wire_13), .Value_2(wire_6), .Written(wire_19));
  mand # (.UUID(64'd1207172339067544539 ^ UUID)) mand_92 (.clk(clk), .rst(rst), .Input_1(wire_34), .Input_2(wire_17), .Output(wire_7));
  mand # (.UUID(64'd1055636189021926738 ^ UUID)) mand_93 (.clk(clk), .rst(rst), .Input_1(wire_16), .Input_2(wire_17), .Output(wire_26));
  mand # (.UUID(64'd3603338431621519469 ^ UUID)) mand_94 (.clk(clk), .rst(rst), .Input_1(wire_37), .Input_2(wire_17), .Output(wire_49));
  OnOrOff # (.UUID(64'd2326604957341175433 ^ UUID)) OnOrOff_95 (.clk(clk), .rst(rst), .Input(wire_18), .Output(wire_17_1));
  TC_Counter # (.UUID(64'd3781882184507484018 ^ UUID), .BIT_WIDTH(64'd64), .count(64'd1)) Counter64_96 (.clk(clk), .rst(rst), .save(wire_39), .in(wire_21), .out(wire_21));

  wire [63:0] wire_0;
  wire [63:0] wire_0_0;
  wire [63:0] wire_0_1;
  wire [63:0] wire_0_2;
  wire [63:0] wire_0_3;
  wire [63:0] wire_0_4;
  wire [63:0] wire_0_5;
  assign wire_0 = wire_0_0|wire_0_1|wire_0_2|wire_0_3|wire_0_4|wire_0_5;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [63:0] wire_4;
  wire [63:0] wire_5;
  wire [63:0] wire_5_0;
  wire [63:0] wire_5_1;
  assign wire_5 = wire_5_0|wire_5_1;
  wire [63:0] wire_6;
  wire [0:0] wire_7;
  wire [63:0] wire_8;
  wire [63:0] wire_8_0;
  wire [63:0] wire_8_1;
  wire [63:0] wire_8_2;
  wire [63:0] wire_8_3;
  assign wire_8 = wire_8_0|wire_8_1|wire_8_2|wire_8_3;
  wire [0:0] wire_9;
  wire [63:0] wire_10;
  wire [63:0] wire_11;
  wire [63:0] wire_12;
  wire [63:0] wire_13;
  wire [63:0] wire_14;
  wire [63:0] wire_14_0;
  wire [63:0] wire_14_1;
  assign wire_14 = wire_14_0|wire_14_1;
  wire [63:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_17_0;
  wire [0:0] wire_17_1;
  wire [0:0] wire_17_2;
  assign wire_17 = wire_17_0|wire_17_1|wire_17_2;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [63:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [63:0] wire_24;
  wire [7:0] wire_25;
  wire [0:0] wire_26;
  wire [63:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [63:0] wire_31;
  wire [0:0] wire_32;
  wire [63:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [7:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_38_0;
  wire [0:0] wire_38_1;
  assign wire_38 = wire_38_0|wire_38_1;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [63:0] wire_42;
  wire [0:0] wire_43;
  wire [63:0] wire_44;
  wire [63:0] wire_45;
  wire [0:0] wire_46;
  wire [63:0] wire_47;
  wire [63:0] wire_48;
  wire [0:0] wire_49;
  wire [63:0] wire_50;
  wire [63:0] wire_50_0;
  wire [63:0] wire_50_1;
  assign wire_50 = wire_50_0|wire_50_1;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_52_0;
  wire [0:0] wire_52_1;
  assign wire_52 = wire_52_0|wire_52_1;
  wire [63:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [0:0] wire_58;
  wire [63:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [63:0] wire_62;
  wire [0:0] wire_63;
  assign wire_63 = 0;
  wire [63:0] wire_64;
  wire [63:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [63:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [63:0] wire_72;
  wire [63:0] wire_73;

endmodule
