module Day3Part2 (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_FileLoader # (.UUID(64'd670867910265240022 ^ UUID), .DEFAULT_FILE_NAME("day3")) FileLoader_0 (.clk(clk), .rst(rst), .en(wire_24), .address(wire_28), .out(wire_17_0));
  TC_Constant # (.UUID(64'd3936697611034503221 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_1 (.out(wire_24));
  TC_FileLoader # (.UUID(64'd1471818332144234541 ^ UUID), .DEFAULT_FILE_NAME("day3_test_1")) FileLoader_2 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_28), .out(wire_17_1));
  TC_Constant # (.UUID(64'd3499631194368056916 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_3 (.out());
  TC_Constant # (.UUID(64'd2232736622141656856 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_4 (.out());
  TC_Constant # (.UUID(64'd1981730186504267880 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_5 (.out());
  TC_Constant # (.UUID(64'd1021525384996764303 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_6 (.out());
  TC_Constant # (.UUID(64'd2233006607170672073 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_7 (.out());
  TC_Constant # (.UUID(64'd2545521340778047509 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_8 (.out());
  TC_Constant # (.UUID(64'd106938163112223798 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_9 (.out());
  TC_Constant # (.UUID(64'd4318802647083067959 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_10 (.out());
  TC_Constant # (.UUID(64'd1130820721428926793 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_11 (.out());
  TC_Constant # (.UUID(64'd291644535782022576 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_12 (.out());
  TC_Constant # (.UUID(64'd4226570772319391860 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_13 (.out());
  TC_Constant # (.UUID(64'd2621130069460615979 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_14 (.out());
  TC_Constant # (.UUID(64'd810286633950345646 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_15 (.out());
  TC_Constant # (.UUID(64'd154484762821244521 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_16 (.out());
  TC_Constant # (.UUID(64'd1293101044721837465 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_17 (.out());
  TC_Constant # (.UUID(64'd1919304839526120989 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFFFFFFFFFFFFFFFF)) Constant64_18 (.out(wire_59));
  TC_Add # (.UUID(64'd539826787227496491 ^ UUID), .BIT_WIDTH(64'd64)) Add64_19 (.in0(wire_61), .in1(wire_20), .ci(1'd0), .out(wire_15), .co());
  TC_DelayLine # (.UUID(64'd1121378025258459254 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_20 (.clk(clk), .rst(rst), .in(wire_15), .out(wire_20));
  TC_Mux # (.UUID(64'd400526689135511509 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_21 (.sel(wire_4), .in0(wire_59), .in1(wire_20), .out(wire_28));
  TC_Switch # (.UUID(64'd3750085722990771933 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_22 (.en(wire_4), .in({{56{1'b0}}, wire_66 }), .out(wire_61));
  TC_Equal # (.UUID(64'd1006503156420949217 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_23 (.in0(wire_20), .in1(wire_37), .out(wire_62));
  TC_And3 # (.UUID(64'd330147788875224171 ^ UUID), .BIT_WIDTH(64'd1)) And3_24 (.in0(wire_56), .in1(wire_36), .in2(wire_74), .out(wire_4));
  TC_Not # (.UUID(64'd285764211932754545 ^ UUID), .BIT_WIDTH(64'd1)) Not_25 (.in(wire_62), .out(wire_74));
  TC_Ram # (.UUID(64'd889594913348838705 ^ UUID), .WORD_WIDTH(64'd128), .WORD_COUNT(64'd512)) Ram_26 (.clk(clk), .rst(rst), .load(wire_18[0:0]), .save(wire_11), .address(wire_0), .in0(wire_44), .in1(wire_41), .in2(64'd0), .in3(64'd0), .out0(wire_12), .out1(wire_19), .out2(), .out3());
  TC_Not # (.UUID(64'd3539672329771887091 ^ UUID), .BIT_WIDTH(64'd1)) Not_27 (.in(wire_5), .out(wire_25));
  TC_Mux # (.UUID(64'd869346753072203086 ^ UUID), .BIT_WIDTH(64'd32)) Mux32_28 (.sel(wire_33), .in0(wire_0), .in1(32'd0), .out(wire_76));
  TC_Not # (.UUID(64'd1498694609800071896 ^ UUID), .BIT_WIDTH(64'd1)) Not_29 (.in(wire_70), .out(wire_23));
  TC_Not # (.UUID(64'd1524827408234024151 ^ UUID), .BIT_WIDTH(64'd1)) Not_30 (.in(wire_53), .out(wire_11));
  TC_And3 # (.UUID(64'd3042879754477079505 ^ UUID), .BIT_WIDTH(64'd1)) And3_31 (.in0(wire_25), .in1(wire_51), .in2(wire_55), .out(wire_70));
  TC_Equal # (.UUID(64'd3161989386235867289 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_32 (.in0(wire_0), .in1(wire_31[31:0]), .out(wire_64));
  TC_Switch # (.UUID(64'd948381973252070923 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_33 (.en(wire_5), .in(wire_0), .out(wire_3));
  TC_Not # (.UUID(64'd1674548457943997484 ^ UUID), .BIT_WIDTH(64'd1)) Not_34 (.in(wire_27), .out(wire_55));
  TC_And # (.UUID(64'd2893488111660484409 ^ UUID), .BIT_WIDTH(64'd1)) And_35 (.in0(wire_64), .in1(wire_50), .out(wire_27));
  TC_Halt # (.UUID(64'd1474802306642119463 ^ UUID), .HALT_MESSAGE("End of file reached!")) Halt_36 (.clk(clk), .rst(rst), .en(wire_52));
  TC_Halt # (.UUID(64'd3727559317572521050 ^ UUID), .HALT_MESSAGE("Found crossing")) Halt_37 (.clk(clk), .rst(rst), .en(1'd0));
  TC_And3 # (.UUID(64'd3134744527415087055 ^ UUID), .BIT_WIDTH(64'd1)) And3_38 (.in0(wire_36), .in1(wire_27), .in2(wire_62), .out(wire_52));
  TC_FileLoader # (.UUID(64'd3429124062269983960 ^ UUID), .DEFAULT_FILE_NAME("day3_test_2")) FileLoader_39 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_28), .out(wire_17_2));
  TC_FileLoader # (.UUID(64'd1473616339079632962 ^ UUID), .DEFAULT_FILE_NAME("day3_test_3")) FileLoader_40 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_28), .out(wire_17_3));
  TC_Halt # (.UUID(64'd2886596719389344914 ^ UUID), .HALT_MESSAGE("Adder overflow! (PositionAdder)")) Halt_41 (.clk(clk), .rst(rst), .en(1'd0));
  TC_DelayLine # (.UUID(64'd4084865240337909835 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_42 (.clk(clk), .rst(rst), .in(wire_44), .out(wire_29));
  TC_Counter # (.UUID(64'd1078548748747073918 ^ UUID), .BIT_WIDTH(64'd32), .count(32'd1)) Counter32_43 (.clk(clk), .rst(rst), .save(wire_33), .in(wire_76), .out(wire_0));
  TC_DelayLine # (.UUID(64'd1099126945014138228 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_44 (.clk(clk), .rst(rst), .in(wire_12), .out(wire_32));
  TC_FileLoader # (.UUID(64'd784893077974596701 ^ UUID), .DEFAULT_FILE_NAME("day3_test_4")) FileLoader_45 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_28), .out(wire_17_4));
  TC_FileLoader # (.UUID(64'd224237426130976828 ^ UUID), .DEFAULT_FILE_NAME("day3_test_5")) FileLoader_46 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_28), .out(wire_17_5));
  TC_FileLoader # (.UUID(64'd4283039450414421346 ^ UUID), .DEFAULT_FILE_NAME("day3_test_6")) FileLoader_47 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_28), .out(wire_17_6));
  TC_FileLoader # (.UUID(64'd1657938444342303651 ^ UUID), .DEFAULT_FILE_NAME("day3_test_7")) FileLoader_48 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_28), .out(wire_17_7));
  TC_NoteSound # (.UUID(64'd428366861129437171 ^ UUID)) NoteSound_49 (.clk(clk), .rst(rst), .command({{7{1'b0}}, wire_52 }), .note(8'd0), .pitch(8'd0));
  TC_Switch # (.UUID(64'd2241906331493591448 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_50 (.en(wire_4), .in(wire_17), .out(wire_60));
  TC_Add # (.UUID(64'd3720721045896377580 ^ UUID), .BIT_WIDTH(64'd64)) Add64_51 (.in0(wire_30), .in1({{48{1'b0}}, wire_21 }), .ci(1'd0), .out(wire_41), .co());
  TC_DelayLine # (.UUID(64'd35903268895255636 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_52 (.clk(clk), .rst(rst), .in(wire_41), .out(wire_30));
  TC_Splitter32 # (.UUID(64'd4160806008740110644 ^ UUID)) Splitter32_53 (.in(wire_14), .out0(wire_63), .out1(wire_73), .out2(), .out3());
  TC_Maker16 # (.UUID(64'd2298888647381191589 ^ UUID)) Maker16_54 (.in0(wire_63), .in1(wire_73), .out(wire_21));
  TC_Splitter32 # (.UUID(64'd3575585577948491953 ^ UUID)) Splitter32_55 (.in(wire_14), .out0(wire_57), .out1(wire_38), .out2(), .out3());
  TC_Maker16 # (.UUID(64'd2926696989604587844 ^ UUID)) Maker16_56 (.in0(wire_57), .in1(wire_38), .out(wire_67));
  TC_Mux # (.UUID(64'd3613559239380446680 ^ UUID), .BIT_WIDTH(64'd32)) Mux32_57 (.sel(wire_49), .in0(wire_58), .in1(wire_7), .out(wire_47));
  TC_DelayLine # (.UUID(64'd1602588821381884070 ^ UUID), .BIT_WIDTH(64'd32)) DelayLine32_58 (.clk(clk), .rst(rst), .in(wire_47), .out(wire_7));
  TC_Add # (.UUID(64'd814287441108641455 ^ UUID), .BIT_WIDTH(64'd32)) Add32_59 (.in0({{16{1'b0}}, wire_67 }), .in1(wire_7), .ci(1'd0), .out(wire_58), .co());
  TC_Not # (.UUID(64'd1441814802550084725 ^ UUID), .BIT_WIDTH(64'd1)) Not_60 (.in(wire_27), .out(wire_49));
  TC_Add # (.UUID(64'd3994601476181792906 ^ UUID), .BIT_WIDTH(64'd32)) Add32_61 (.in0(wire_19[31:0]), .in1(wire_47), .ci(1'd0), .out(wire_9), .co());
  TC_Add # (.UUID(64'd1265684793700429268 ^ UUID), .BIT_WIDTH(64'd32)) Add32_62 (.in0(wire_9), .in1(wire_26), .ci(1'd0), .out(wire_43), .co());
  TC_Switch # (.UUID(64'd474332149679910780 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_63 (.en(wire_45), .in(wire_43), .out(wire_54));
  InputMananger # (.UUID(64'd280349663464583758 ^ UUID)) InputMananger_64 (.clk(clk), .rst(rst), .Main_8b(wire_60), .Offset(wire_66), .Output(wire_14), .NewLine(wire_5));
  QuickSave # (.UUID(64'd3964331221245691836 ^ UUID)) QuickSave_65 (.clk(clk), .rst(rst), .Value(wire_17), .\Number_(stored) (wire_37), .\Saved?_1 (wire_36), .\Saved?_2 (wire_51));
  ManhattanDistance # (.UUID(64'd4534475870914388036 ^ UUID)) ManhattanDistance_66 (.clk(clk), .rst(rst), .X(wire_40), .Y(wire_72), .Output(wire_65));
  CellRotator # (.UUID(64'd2988738449177159528 ^ UUID)) CellRotator_67 (.clk(clk), .rst(rst), .Tick(wire_27), .Input(wire_39), .Pos_2(wire_13), .Pos_1(wire_46), .Written());
  QuickSave # (.UUID(64'd3551179199781681902 ^ UUID)) QuickSave_68 (.clk(clk), .rst(rst), .Value({{63{1'b0}}, wire_5 }), .\Number_(stored) (wire_18), .\Saved?_1 (wire_53), .\Saved?_2 ());
  OnOrOff # (.UUID(64'd2880407376120648954 ^ UUID)) OnOrOff_69 (.clk(clk), .rst(rst), .Input(wire_23), .Output(wire_33));
  QuickSave # (.UUID(64'd4013860832325939171 ^ UUID)) QuickSave_70 (.clk(clk), .rst(rst), .Value({{32{1'b0}}, wire_3 }), .\Number_(stored) (wire_31), .\Saved?_1 (wire_50), .\Saved?_2 ());
  OnOrOff # (.UUID(64'd685402883028759750 ^ UUID)) OnOrOff_71 (.clk(clk), .rst(rst), .Input(wire_11), .Output(wire_56_0));
  OnOrOff # (.UUID(64'd2586521289870388092 ^ UUID)) OnOrOff_72 (.clk(clk), .rst(rst), .Input(wire_27), .Output(wire_56_1));
  PositionAdder # (.UUID(64'd1952379698983790479 ^ UUID)) PositionAdder_73 (.clk(clk), .rst(rst), .Current_Position(wire_29), .Move({{32{1'b0}}, wire_14 }), .overflow(wire_75), .New_Position(wire_44));
  PositionAdder # (.UUID(64'd549660374295142354 ^ UUID)) PositionAdder_74 (.clk(clk), .rst(rst), .Current_Position(wire_13), .Move({{32{1'b0}}, wire_14 }), .overflow(), .New_Position(wire_39));
  LineCrosserz_3 # (.UUID(64'd235678000759494782 ^ UUID)) LineCrosserz_3_75 (.clk(clk), .rst(rst), .L2End(wire_13), .L2Start(wire_46), .L1End(wire_12), .L1Start(wire_32), .Intercection(wire_45), .Point_of_Interce(wire_2), .\StepCount_(r) (wire_16));
  _64bz_toz_32b # (.UUID(64'd4074607966076726035 ^ UUID)) _64bz_toz_32b_76 (.clk(clk), .rst(rst), .Input(wire_32), .Output_1(wire_35), .Output_2(wire_34));
  _64bz_toz_32b # (.UUID(64'd3297953936306396081 ^ UUID)) _64bz_toz_32b_77 (.clk(clk), .rst(rst), .Input(wire_12), .Output_1(wire_42), .Output_2(wire_22));
  _64bz_toz_32b # (.UUID(64'd2799350786039608227 ^ UUID)) _64bz_toz_32b_78 (.clk(clk), .rst(rst), .Input(wire_46), .Output_1(wire_68), .Output_2(wire_1));
  _64bz_toz_32b # (.UUID(64'd4547022319690718172 ^ UUID)) _64bz_toz_32b_79 (.clk(clk), .rst(rst), .Input(wire_13), .Output_1(wire_10), .Output_2(wire_6));
  _64bz_toz_32b # (.UUID(64'd36584691338760372 ^ UUID)) _64bz_toz_32b_80 (.clk(clk), .rst(rst), .Input(wire_2), .Output_1(wire_72), .Output_2(wire_40));
  _64bz_toz_32b # (.UUID(64'd1683694981542803589 ^ UUID)) _64bz_toz_32b_81 (.clk(clk), .rst(rst), .Input(wire_29), .Output_1(wire_69), .Output_2(wire_8));
  NumberDisplayz_zmz_1rzm10d # (.UUID(64'd1558355514723882557 ^ UUID)) NumberDisplayz_zmz_1rzm10d_82 (.clk(clk), .rst(rst), .Input(wire_8));
  NumberDisplayz_zmz_1rzm10d # (.UUID(64'd1342504794432391415 ^ UUID)) NumberDisplayz_zmz_1rzm10d_83 (.clk(clk), .rst(rst), .Input(wire_69));
  Minimuum # (.UUID(64'd1847184604891007288 ^ UUID)) Minimuum_84 (.clk(clk), .rst(rst), .Value({{32{1'b0}}, wire_54 }), .Smallest(wire_71));
  NumberDisplayz_zmz_1rzm10d # (.UUID(64'd17818789641386411 ^ UUID)) NumberDisplayz_zmz_1rzm10d_85 (.clk(clk), .rst(rst), .Input(wire_71[31:0]));
  Minimuum # (.UUID(64'd3754522689005736836 ^ UUID)) Minimuum_86 (.clk(clk), .rst(rst), .Value({{32{1'b0}}, wire_65 }), .Smallest(wire_48));
  NumberDisplayz_zmz_1rzm10d # (.UUID(64'd3168566118355095045 ^ UUID)) NumberDisplayz_zmz_1rzm10d_87 (.clk(clk), .rst(rst), .Input(wire_48[31:0]));
  InverseAbs32b # (.UUID(64'd1716325306459498110 ^ UUID)) InverseAbs32b_88 (.clk(clk), .rst(rst), .Input(wire_16), .Output(wire_26));

  wire [31:0] wire_0;
  wire [31:0] wire_1;
  wire [63:0] wire_2;
  wire [31:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [31:0] wire_6;
  wire [31:0] wire_7;
  wire [31:0] wire_8;
  wire [31:0] wire_9;
  wire [31:0] wire_10;
  wire [0:0] wire_11;
  wire [63:0] wire_12;
  wire [63:0] wire_13;
  wire [31:0] wire_14;
  wire [63:0] wire_15;
  wire [31:0] wire_16;
  wire [63:0] wire_17;
  wire [63:0] wire_17_0;
  wire [63:0] wire_17_1;
  wire [63:0] wire_17_2;
  wire [63:0] wire_17_3;
  wire [63:0] wire_17_4;
  wire [63:0] wire_17_5;
  wire [63:0] wire_17_6;
  wire [63:0] wire_17_7;
  assign wire_17 = wire_17_0|wire_17_1|wire_17_2|wire_17_3|wire_17_4|wire_17_5|wire_17_6|wire_17_7;
  wire [63:0] wire_18;
  wire [63:0] wire_19;
  wire [63:0] wire_20;
  wire [15:0] wire_21;
  wire [31:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [31:0] wire_26;
  wire [0:0] wire_27;
  wire [63:0] wire_28;
  wire [63:0] wire_29;
  wire [63:0] wire_30;
  wire [63:0] wire_31;
  wire [63:0] wire_32;
  wire [0:0] wire_33;
  wire [31:0] wire_34;
  wire [31:0] wire_35;
  wire [0:0] wire_36;
  wire [63:0] wire_37;
  wire [7:0] wire_38;
  wire [63:0] wire_39;
  wire [31:0] wire_40;
  wire [63:0] wire_41;
  wire [31:0] wire_42;
  wire [31:0] wire_43;
  wire [63:0] wire_44;
  wire [0:0] wire_45;
  wire [63:0] wire_46;
  wire [31:0] wire_47;
  wire [63:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [31:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_56_0;
  wire [0:0] wire_56_1;
  assign wire_56 = wire_56_0|wire_56_1;
  wire [7:0] wire_57;
  wire [31:0] wire_58;
  wire [63:0] wire_59;
  wire [63:0] wire_60;
  wire [63:0] wire_61;
  wire [0:0] wire_62;
  wire [7:0] wire_63;
  wire [0:0] wire_64;
  wire [31:0] wire_65;
  wire [7:0] wire_66;
  wire [15:0] wire_67;
  wire [31:0] wire_68;
  wire [31:0] wire_69;
  wire [0:0] wire_70;
  wire [63:0] wire_71;
  wire [31:0] wire_72;
  wire [7:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [31:0] wire_76;

endmodule
