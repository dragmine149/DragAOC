module InputMananger (clk, rst, Main_8b, Offset, Output, NewLine);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [63:0] Main_8b;
  output  wire [7:0] Offset;
  output  wire [31:0] Output;
  output  wire [0:0] NewLine;

  TC_Not # (.UUID(64'd931508675602096990 ^ UUID), .BIT_WIDTH(64'd1)) Not_0 (.in(wire_35), .out(wire_8));
  TC_Not # (.UUID(64'd3022390878210203468 ^ UUID), .BIT_WIDTH(64'd1)) Not_1 (.in(wire_14), .out(wire_40));
  TC_Not # (.UUID(64'd1800283864298422345 ^ UUID), .BIT_WIDTH(64'd1)) Not_2 (.in(wire_26), .out(wire_18));
  TC_IndexerByte # (.UUID(64'd97685308338425177 ^ UUID), .INDEX(64'd0)) IndexerByte_3 (.in(wire_20), .out(wire_43));
  TC_IndexerByte # (.UUID(64'd1535575929618738446 ^ UUID), .INDEX(64'd1)) IndexerByte_4 (.in(wire_20), .out(wire_4));
  TC_IndexerByte # (.UUID(64'd2193632466719870419 ^ UUID), .INDEX(64'd2)) IndexerByte_5 (.in(wire_20), .out(wire_11));
  TC_IndexerByte # (.UUID(64'd2107427035108924588 ^ UUID), .INDEX(64'd3)) IndexerByte_6 (.in(wire_20), .out(wire_41));
  TC_IndexerByte # (.UUID(64'd3440309831824146801 ^ UUID), .INDEX(64'd4)) IndexerByte_7 (.in(wire_20), .out(wire_17));
  TC_Not # (.UUID(64'd3291242525983120137 ^ UUID), .BIT_WIDTH(64'd1)) Not_8 (.in(wire_42), .out(wire_22));
  TC_Not # (.UUID(64'd3621447621843358213 ^ UUID), .BIT_WIDTH(64'd1)) Not_9 (.in(wire_33), .out(wire_25));
  TC_Constant # (.UUID(64'd4128177160354142202 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_10 (.out(wire_23));
  TC_Constant # (.UUID(64'd1450032060031438387 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_11 (.out(wire_13));
  TC_Constant # (.UUID(64'd720295887030816158 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5)) Constant8_12 (.out(wire_29));
  TC_Switch # (.UUID(64'd1796095839427953768 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_13 (.en(wire_14), .in(wire_12), .out(wire_30));
  TC_Switch # (.UUID(64'd2922149858396693218 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_14 (.en(wire_35), .in(wire_15), .out(wire_27));
  TC_Switch # (.UUID(64'd3922512512722123755 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_15 (.en(wire_8), .in(wire_15), .out(wire_7_3));
  TC_Switch # (.UUID(64'd1661399743869514783 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_16 (.en(wire_16), .in(wire_12), .out(wire_7_2));
  TC_Switch # (.UUID(64'd101279653130619089 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_17 (.en(wire_3), .in(wire_36), .out(wire_7_1));
  TC_Equal # (.UUID(64'd574040698186393 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_18 (.in0(wire_5), .in1(wire_31), .out(wire_21));
  TC_Constant # (.UUID(64'd3169959144025133120 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hA)) Constant8_19 (.out(wire_31));
  TC_Constant # (.UUID(64'd1774062521881063346 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_20 (.out());
  TC_Switch # (.UUID(64'd1663735972669831967 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_21 (.en(wire_8), .in(wire_32), .out(wire_5_3));
  TC_Switch # (.UUID(64'd1682384720783853639 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_22 (.en(wire_16), .in(wire_19), .out(wire_5_2));
  TC_Switch # (.UUID(64'd336630731137340894 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_23 (.en(wire_3), .in(wire_6), .out(wire_5_1));
  TC_Switch # (.UUID(64'd1090600476240894467 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_24 (.en(wire_2), .in(wire_36), .out(wire_7_0));
  TC_Constant # (.UUID(64'd1929537234046566558 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_25 (.out(wire_10));
  TC_IndexerByte # (.UUID(64'd4141135529995031329 ^ UUID), .INDEX(64'd5)) IndexerByte_26 (.in(wire_20), .out(wire_34));
  ByteToNumbersz_2 # (.UUID(64'd4133949311826805421 ^ UUID)) ByteToNumbersz_2_27 (.clk(clk), .rst(rst), .Input(wire_17), .Has_48(wire_26), .Number(wire_6));
  ByteToNumbersz_2 # (.UUID(64'd1272090532466054217 ^ UUID)) ByteToNumbersz_2_28 (.clk(clk), .rst(rst), .Input(wire_41), .Has_48(wire_14), .Number(wire_19));
  ByteToNumbersz_2 # (.UUID(64'd442016588560264049 ^ UUID)) ByteToNumbersz_2_29 (.clk(clk), .rst(rst), .Input(wire_11), .Has_48(wire_35), .Number(wire_32));
  ByteToNumbersz_2 # (.UUID(64'd2890634684432758681 ^ UUID)) ByteToNumbersz_2_30 (.clk(clk), .rst(rst), .Input(wire_4), .Has_48(), .Number(wire_39));
  OnOrOff # (.UUID(64'd1293384845730880674 ^ UUID)) OnOrOff_31 (.clk(clk), .rst(rst), .Input(wire_8), .Output(wire_42));
  OnOrOff # (.UUID(64'd1199503870914616836 ^ UUID)) OnOrOff_32 (.clk(clk), .rst(rst), .Input(wire_42), .Output(wire_33_1));
  mand # (.UUID(64'd71773308005596248 ^ UUID)) mand_33 (.clk(clk), .rst(rst), .Input_1(wire_22), .Input_2(wire_40), .Output(wire_16));
  OnOrOff # (.UUID(64'd2496479277812182200 ^ UUID)) OnOrOff_34 (.clk(clk), .rst(rst), .Input(wire_16), .Output(wire_33_0));
  OnOrOff # (.UUID(64'd562383047764755250 ^ UUID)) OnOrOff_35 (.clk(clk), .rst(rst), .Input(wire_33), .Output(wire_1_0));
  mand # (.UUID(64'd2207443847502782851 ^ UUID)) mand_36 (.clk(clk), .rst(rst), .Input_1(wire_25), .Input_2(wire_18), .Output(wire_3));
  OnOrOff # (.UUID(64'd4599396002788419685 ^ UUID)) OnOrOff_37 (.clk(clk), .rst(rst), .Input(wire_3), .Output(wire_1_1));
  _8rSwitch # (.UUID(64'd1575133784720396750 ^ UUID)) _8rSwitch_38 (.clk(clk), .rst(rst), .Enable(wire_8), .Input(wire_23), .Output(wire_0_3));
  _8rSwitch # (.UUID(64'd4543931877293036313 ^ UUID)) _8rSwitch_39 (.clk(clk), .rst(rst), .Enable(wire_16), .Input(wire_13), .Output(wire_0_2));
  _8rSwitch # (.UUID(64'd1095850944845713730 ^ UUID)) _8rSwitch_40 (.clk(clk), .rst(rst), .Enable(wire_3), .Input(wire_29), .Output(wire_0_1));
  ByteToDirection # (.UUID(64'd2513996509828058476 ^ UUID)) ByteToDirection_41 (.clk(clk), .rst(rst), .Input(wire_43), .Bit_1(wire_37), .Bit_2(wire_24));
  x10zpnz_ZL16bZR # (.UUID(64'd723796272159468420 ^ UUID)) x10zpnz_ZL16bZR_42 (.clk(clk), .rst(rst), .Input_1(wire_19), .Input_2(wire_27), .Output(wire_12));
  x10zpnz_ZL16bZR # (.UUID(64'd1036033709405592105 ^ UUID)) x10zpnz_ZL16bZR_43 (.clk(clk), .rst(rst), .Input_1(wire_32), .Input_2({{8{1'b0}}, wire_39 }), .Output(wire_15));
  x10zpnz_ZL16bZR # (.UUID(64'd3635845447600608103 ^ UUID)) x10zpnz_ZL16bZR_44 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_30), .Output(wire_36));
  Translator # (.UUID(64'd615318436903473277 ^ UUID)) Translator_45 (.clk(clk), .rst(rst), .Input_1(wire_7), .Input_2(wire_37), .Input_3(wire_24), .Output(wire_28));
  _8rSwitch # (.UUID(64'd3085616695338917016 ^ UUID)) _8rSwitch_46 (.clk(clk), .rst(rst), .Enable(wire_2), .Input(wire_10), .Output(wire_0_0));
  ByteToNumbersz_2 # (.UUID(64'd2537531887911040497 ^ UUID)) ByteToNumbersz_2_47 (.clk(clk), .rst(rst), .Input(wire_34), .Has_48(), .Number(wire_38));
  _8rSwitch # (.UUID(64'd42025438754252433 ^ UUID)) _8rSwitch_48 (.clk(clk), .rst(rst), .Enable(wire_2), .Input(wire_38), .Output(wire_5_0));
  mand # (.UUID(64'd1787362092892007500 ^ UUID)) mand_49 (.clk(clk), .rst(rst), .Input_1(wire_26), .Input_2(wire_9), .Output(wire_2));
  TC_Not # (.UUID(64'd48304628449859450 ^ UUID), .BIT_WIDTH(64'd1)) Not_50 (.in(wire_1), .out(wire_9));

  wire [7:0] wire_0;
  wire [7:0] wire_0_0;
  wire [7:0] wire_0_1;
  wire [7:0] wire_0_2;
  wire [7:0] wire_0_3;
  assign wire_0 = wire_0_0|wire_0_1|wire_0_2|wire_0_3;
  assign Offset = wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_1_0;
  wire [0:0] wire_1_1;
  assign wire_1 = wire_1_0|wire_1_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  wire [7:0] wire_5;
  wire [7:0] wire_5_0;
  wire [7:0] wire_5_1;
  wire [7:0] wire_5_2;
  wire [7:0] wire_5_3;
  assign wire_5 = wire_5_0|wire_5_1|wire_5_2|wire_5_3;
  wire [7:0] wire_6;
  wire [15:0] wire_7;
  wire [15:0] wire_7_0;
  wire [15:0] wire_7_1;
  wire [15:0] wire_7_2;
  wire [15:0] wire_7_3;
  assign wire_7 = wire_7_0|wire_7_1|wire_7_2|wire_7_3;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [7:0] wire_11;
  wire [15:0] wire_12;
  wire [7:0] wire_13;
  wire [0:0] wire_14;
  wire [15:0] wire_15;
  wire [0:0] wire_16;
  wire [7:0] wire_17;
  wire [0:0] wire_18;
  wire [7:0] wire_19;
  wire [63:0] wire_20;
  assign wire_20 = Main_8b;
  wire [0:0] wire_21;
  assign NewLine = wire_21;
  wire [0:0] wire_22;
  wire [7:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [15:0] wire_27;
  wire [31:0] wire_28;
  assign Output = wire_28;
  wire [7:0] wire_29;
  wire [15:0] wire_30;
  wire [7:0] wire_31;
  wire [7:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_33_0;
  wire [0:0] wire_33_1;
  assign wire_33 = wire_33_0|wire_33_1;
  wire [7:0] wire_34;
  wire [0:0] wire_35;
  wire [15:0] wire_36;
  wire [0:0] wire_37;
  wire [7:0] wire_38;
  wire [7:0] wire_39;
  wire [0:0] wire_40;
  wire [7:0] wire_41;
  wire [0:0] wire_42;
  wire [7:0] wire_43;

endmodule
