module LineCrosserz_3 (clk, rst, Input_1, Input_2, Input_3, Input_4, Output_1, Output_2);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [31:0] Input_1;
  input  wire [31:0] Input_2;
  input  wire [31:0] Input_3;
  input  wire [31:0] Input_4;
  output  wire [0:0] Output_1;
  output  wire [31:0] Output_2;

  TC_Equal # (.UUID(64'd4270302367443503270 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_0 (.in0(wire_38), .in1(wire_50), .out(wire_10));
  TC_Equal # (.UUID(64'd610006227766373642 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_1 (.in0(wire_21), .in1(wire_27), .out(wire_46));
  TC_Equal # (.UUID(64'd115549839275673676 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_2 (.in0(wire_35), .in1(wire_37), .out(wire_9));
  TC_Equal # (.UUID(64'd2107797086179499841 ^ UUID), .BIT_WIDTH(64'd16)) Equal16_3 (.in0(wire_28), .in1(wire_5), .out(wire_7));
  TC_Switch # (.UUID(64'd2832402715206588669 ^ UUID), .BIT_WIDTH(64'd32)) Output32z_4 (.en(wire_36), .in(wire_42), .out(Output_2));
  TC_Switch # (.UUID(64'd29451040430517838 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_5 (.en(wire_32), .in(wire_4), .out(wire_23));
  TC_Not # (.UUID(64'd380166382871947097 ^ UUID), .BIT_WIDTH(64'd1)) Not_6 (.in(wire_11), .out(wire_32));
  TC_Switch # (.UUID(64'd1168352118892452644 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_7 (.en(wire_23), .in(wire_18), .out(wire_25_1));
  TC_Switch # (.UUID(64'd3818630122358164471 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_8 (.en(wire_6), .in(wire_18), .out(wire_2_1));
  TC_Switch # (.UUID(64'd371305226280118364 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_9 (.en(wire_6), .in(wire_12), .out(wire_25_0));
  TC_Switch # (.UUID(64'd4219178858152753453 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_10 (.en(wire_23), .in(wire_12), .out(wire_2_0));
  TC_Switch # (.UUID(64'd3821448631046911694 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_11 (.en(wire_43), .in(wire_11), .out(wire_6));
  TC_Not # (.UUID(64'd569669821514979918 ^ UUID), .BIT_WIDTH(64'd1)) Not_12 (.in(wire_23), .out(wire_43));
  TC_Splitter16 # (.UUID(64'd3797087622397082436 ^ UUID)) Splitter16_13 (.in(wire_14), .out0(wire_54), .out1(wire_34));
  TC_Splitter16 # (.UUID(64'd2392608650595757673 ^ UUID)) Splitter16_14 (.in(wire_0), .out0(wire_55), .out1(wire_39));
  TC_Maker32 # (.UUID(64'd16555111681801296 ^ UUID)) Maker32_15 (.in0(wire_55), .in1(wire_39), .in2(wire_54), .in3(wire_34), .out(wire_42));
  TC_And3 # (.UUID(64'd1658388512215494880 ^ UUID), .BIT_WIDTH(64'd1)) And3_16 (.in0(wire_48), .in1(wire_51), .in2(wire_13), .out(wire_36));
  PositionDecoder # (.UUID(64'd3728414520355176465 ^ UUID)) PositionDecoder_17 (.clk(clk), .rst(rst), .Position(wire_33), .Y(wire_5), .X(wire_37));
  PositionDecoder # (.UUID(64'd3687752940276849781 ^ UUID)) PositionDecoder_18 (.clk(clk), .rst(rst), .Position(wire_30), .Y(wire_28), .X(wire_35));
  PositionDecoder # (.UUID(64'd3226381494125033591 ^ UUID)) PositionDecoder_19 (.clk(clk), .rst(rst), .Position(wire_17), .Y(wire_27), .X(wire_50));
  PositionDecoder # (.UUID(64'd2722932116695844045 ^ UUID)) PositionDecoder_20 (.clk(clk), .rst(rst), .Position(wire_26), .Y(wire_21), .X(wire_38));
  _32bz_toz_64b # (.UUID(64'd3154309438596456414 ^ UUID)) _32bz_toz_64b_21 (.clk(clk), .rst(rst), .Input_1(wire_17), .Input_2(wire_26), .Output(wire_18));
  _32bz_toz_64b # (.UUID(64'd2473331021217161339 ^ UUID)) _32bz_toz_64b_22 (.clk(clk), .rst(rst), .Input_1(wire_33), .Input_2(wire_30), .Output(wire_12));
  _64bToPosition # (.UUID(64'd3110367828946421310 ^ UUID)) _64bToPosition_23 (.clk(clk), .rst(rst), .Input(wire_2), .EndY(wire_47), .EndX(), .StartY(wire_31), .StartX(wire_0));
  _64bToPosition # (.UUID(64'd3971100450210234737 ^ UUID)) _64bToPosition_24 (.clk(clk), .rst(rst), .Input(wire_25), .EndY(), .EndX(wire_19), .StartY(wire_14), .StartX(wire_8));
  minmax # (.UUID(64'd1642526826406692316 ^ UUID)) minmax_25 (.clk(clk), .rst(rst), .Input_1(wire_31), .Input_2(wire_47), .Minimum(wire_1), .Maximum(wire_3));
  mand # (.UUID(64'd3025706981059298082 ^ UUID)) mand_26 (.clk(clk), .rst(rst), .Input_1(wire_29), .Input_2(wire_41), .Output(wire_56));
  mand # (.UUID(64'd3923050422831829113 ^ UUID)) mand_27 (.clk(clk), .rst(rst), .Input_1(wire_22), .Input_2(wire_15), .Output(wire_52));
  mand # (.UUID(64'd3934257394102842263 ^ UUID)) mand_28 (.clk(clk), .rst(rst), .Input_1(wire_52), .Input_2(wire_56), .Output(wire_13));
  mand # (.UUID(64'd1966732459903081054 ^ UUID)) mand_29 (.clk(clk), .rst(rst), .Input_1(wire_10), .Input_2(wire_7), .Output(wire_11));
  mand # (.UUID(64'd1967875822324122093 ^ UUID)) mand_30 (.clk(clk), .rst(rst), .Input_1(wire_46), .Input_2(wire_9), .Output(wire_4));
  gte # (.UUID(64'd1912638743888257692 ^ UUID)) gte_31 (.clk(clk), .rst(rst), .Input_1(wire_1), .Input_2(wire_14), .Output(wire_41));
  lte # (.UUID(64'd4471518355096608102 ^ UUID)) lte_32 (.clk(clk), .rst(rst), .Input_1(wire_3), .Input_2(wire_14), .Output(wire_29));
  gte # (.UUID(64'd2526412827706897184 ^ UUID)) gte_33 (.clk(clk), .rst(rst), .Input_1(wire_45), .Input_2(wire_0), .Output(wire_15));
  lte # (.UUID(64'd4451336207933505359 ^ UUID)) lte_34 (.clk(clk), .rst(rst), .Input_1(wire_49), .Input_2(wire_0), .Output(wire_22));
  mOR # (.UUID(64'd3811154444398219071 ^ UUID)) mOR_35 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_23), .Output(wire_51));
  minmax # (.UUID(64'd3928075902182458356 ^ UUID)) minmax_36 (.clk(clk), .rst(rst), .Input_1(wire_8), .Input_2(wire_19), .Minimum(wire_45), .Maximum(wire_49));
  mand # (.UUID(64'd2282199498514448531 ^ UUID)) mand_37 (.clk(clk), .rst(rst), .Input_1(wire_20), .Input_2(wire_53), .Output(wire_40));
  mand # (.UUID(64'd4236102916636182286 ^ UUID)) mand_38 (.clk(clk), .rst(rst), .Input_1(wire_44), .Input_2(wire_24), .Output(wire_16));
  mNOR # (.UUID(64'd1044973136834131328 ^ UUID)) mNOR_39 (.clk(clk), .rst(rst), .Input_1(wire_16), .Input_2(wire_40), .Output(wire_48));
  is0z_32b # (.UUID(64'd683255215662450355 ^ UUID)) is0z_32b_40 (.clk(clk), .rst(rst), .Input(wire_33), .Output(wire_24));
  is0z_32b # (.UUID(64'd2032268312256396280 ^ UUID)) is0z_32b_41 (.clk(clk), .rst(rst), .Input(wire_30), .Output(wire_44));
  is0z_32b # (.UUID(64'd3014373814176874017 ^ UUID)) is0z_32b_42 (.clk(clk), .rst(rst), .Input(wire_17), .Output(wire_53));
  is0z_32b # (.UUID(64'd2506635687769368550 ^ UUID)) is0z_32b_43 (.clk(clk), .rst(rst), .Input(wire_26), .Output(wire_20));

  wire [15:0] wire_0;
  wire [15:0] wire_1;
  wire [63:0] wire_2;
  wire [63:0] wire_2_0;
  wire [63:0] wire_2_1;
  assign wire_2 = wire_2_0|wire_2_1;
  wire [15:0] wire_3;
  wire [0:0] wire_4;
  wire [15:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [15:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [63:0] wire_12;
  wire [0:0] wire_13;
  wire [15:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [31:0] wire_17;
  assign wire_17 = Input_3;
  wire [63:0] wire_18;
  wire [15:0] wire_19;
  wire [0:0] wire_20;
  wire [15:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [63:0] wire_25;
  wire [63:0] wire_25_0;
  wire [63:0] wire_25_1;
  assign wire_25 = wire_25_0|wire_25_1;
  wire [31:0] wire_26;
  assign wire_26 = Input_4;
  wire [15:0] wire_27;
  wire [15:0] wire_28;
  wire [0:0] wire_29;
  wire [31:0] wire_30;
  assign wire_30 = Input_2;
  wire [15:0] wire_31;
  wire [0:0] wire_32;
  wire [31:0] wire_33;
  assign wire_33 = Input_1;
  wire [7:0] wire_34;
  wire [15:0] wire_35;
  wire [0:0] wire_36;
  assign Output_1 = wire_36;
  wire [15:0] wire_37;
  wire [15:0] wire_38;
  wire [7:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [31:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [15:0] wire_45;
  wire [0:0] wire_46;
  wire [15:0] wire_47;
  wire [0:0] wire_48;
  wire [15:0] wire_49;
  wire [15:0] wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [7:0] wire_54;
  wire [7:0] wire_55;
  wire [0:0] wire_56;

endmodule
