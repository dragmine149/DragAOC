module LineCrosserz_3 (clk, rst, L2End, L2Start, L1End, L1Start, Output_1, Output_2);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [63:0] L2End;
  input  wire [63:0] L2Start;
  input  wire [63:0] L1End;
  input  wire [63:0] L1Start;
  output  wire [0:0] Output_1;
  output  wire [63:0] Output_2;

  TC_Switch # (.UUID(64'd29451040430517838 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_0 (.en(wire_10), .in(wire_36), .out(wire_4));
  TC_Not # (.UUID(64'd380166382871947097 ^ UUID), .BIT_WIDTH(64'd1)) Not_1 (.in(wire_23), .out(wire_10));
  TC_Switch # (.UUID(64'd3821448631046911694 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_2 (.en(wire_11), .in(wire_23), .out(wire_22));
  TC_Not # (.UUID(64'd569669821514979918 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_4), .out(wire_11));
  TC_And3 # (.UUID(64'd1658388512215494880 ^ UUID), .BIT_WIDTH(64'd1)) And3_4 (.in0(wire_14), .in1(wire_33), .in2(wire_31), .out(wire_25));
  TC_Equal # (.UUID(64'd1462953451613577458 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_5 (.in0(wire_3), .in1(wire_5), .out(wire_34));
  TC_Equal # (.UUID(64'd2477445908053147713 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_6 (.in0(wire_2), .in1(wire_20), .out(wire_30));
  TC_Equal # (.UUID(64'd3736993343762613191 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_7 (.in0(wire_13), .in1(wire_29), .out(wire_9));
  TC_Equal # (.UUID(64'd2800749848815207265 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_8 (.in0(wire_26), .in1(wire_21), .out(wire_15));
  TC_Switch # (.UUID(64'd1144186547777792254 ^ UUID), .BIT_WIDTH(64'd64)) Output64z_9 (.en(wire_25), .in(wire_17), .out(Output_2));
  TC_Constant # (.UUID(64'd1651574857256674590 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_10 (.out());
  mand # (.UUID(64'd1966732459903081054 ^ UUID)) mand_11 (.clk(clk), .rst(rst), .Input_1(wire_34), .Input_2(wire_15), .Output(wire_23));
  mand # (.UUID(64'd1967875822324122093 ^ UUID)) mand_12 (.clk(clk), .rst(rst), .Input_1(wire_30), .Input_2(wire_9), .Output(wire_36));
  mOR # (.UUID(64'd3811154444398219071 ^ UUID)) mOR_13 (.clk(clk), .rst(rst), .Input_1(wire_4), .Input_2(wire_22), .Output(wire_33));
  mand # (.UUID(64'd2282199498514448531 ^ UUID)) mand_14 (.clk(clk), .rst(rst), .Input_1(wire_32), .Input_2(wire_12), .Output(wire_35));
  mand # (.UUID(64'd4236102916636182286 ^ UUID)) mand_15 (.clk(clk), .rst(rst), .Input_1(wire_1), .Input_2(wire_19), .Output(wire_27));
  mNOR # (.UUID(64'd1044973136834131328 ^ UUID)) mNOR_16 (.clk(clk), .rst(rst), .Input_1(wire_27), .Input_2(wire_35), .Output(wire_14));
  _64bz_toz_32b # (.UUID(64'd1160700702824551150 ^ UUID)) _64bz_toz_32b_17 (.clk(clk), .rst(rst), .Input(wire_16), .Output_1(wire_21), .Output_2(wire_29));
  _64bz_toz_32b # (.UUID(64'd4249573345702729115 ^ UUID)) _64bz_toz_32b_18 (.clk(clk), .rst(rst), .Input(wire_24), .Output_1(wire_26), .Output_2(wire_13));
  _64bz_toz_32b # (.UUID(64'd3482476773988014960 ^ UUID)) _64bz_toz_32b_19 (.clk(clk), .rst(rst), .Input(wire_0), .Output_1(wire_20), .Output_2(wire_5));
  _64bz_toz_32b # (.UUID(64'd1881820232260440322 ^ UUID)) _64bz_toz_32b_20 (.clk(clk), .rst(rst), .Input(wire_28), .Output_1(wire_2), .Output_2(wire_3));
  is0z_64b # (.UUID(64'd3522606142968185792 ^ UUID)) is0z_64b_21 (.clk(clk), .rst(rst), .Input(wire_28), .Output(wire_32));
  is0z_64b # (.UUID(64'd2383929583881890307 ^ UUID)) is0z_64b_22 (.clk(clk), .rst(rst), .Input(wire_0), .Output(wire_12));
  is0z_64b # (.UUID(64'd3448954266748536719 ^ UUID)) is0z_64b_23 (.clk(clk), .rst(rst), .Input(wire_24), .Output(wire_1));
  is0z_64b # (.UUID(64'd908196902127981698 ^ UUID)) is0z_64b_24 (.clk(clk), .rst(rst), .Input(wire_16), .Output(wire_19));
  PositionChcker # (.UUID(64'd470197739512970021 ^ UUID)) PositionChcker_25 (.clk(clk), .rst(rst), .HorizontalEnd(wire_8), .VerticalEnd(wire_7), .VerticalStart(wire_18), .HorizontalStart(wire_6), .Output_1(wire_31), .Output_2(wire_17));
  BusSwitcher # (.UUID(64'd4508613529556397755 ^ UUID)) BusSwitcher_26 (.clk(clk), .rst(rst), .Line_End(wire_0), .Line_Start(wire_28), .Option_1(wire_22), .Option_2(wire_4), .Horizontal_End(wire_8_1), .Horizontal_Start(wire_6_0), .Vertical_End(wire_7_1), .Vertical_Start(wire_18_0));
  BusSwitcher # (.UUID(64'd1656550384719575395 ^ UUID)) BusSwitcher_27 (.clk(clk), .rst(rst), .Line_End(wire_16), .Line_Start(wire_24), .Option_1(wire_4), .Option_2(wire_22), .Horizontal_End(wire_8_0), .Horizontal_Start(wire_6_1), .Vertical_End(wire_7_0), .Vertical_Start(wire_18_1));

  wire [63:0] wire_0;
  assign wire_0 = L1End;
  wire [0:0] wire_1;
  wire [31:0] wire_2;
  wire [31:0] wire_3;
  wire [0:0] wire_4;
  wire [31:0] wire_5;
  wire [63:0] wire_6;
  wire [63:0] wire_6_0;
  wire [63:0] wire_6_1;
  assign wire_6 = wire_6_0|wire_6_1;
  wire [63:0] wire_7;
  wire [63:0] wire_7_0;
  wire [63:0] wire_7_1;
  assign wire_7 = wire_7_0|wire_7_1;
  wire [63:0] wire_8;
  wire [63:0] wire_8_0;
  wire [63:0] wire_8_1;
  assign wire_8 = wire_8_0|wire_8_1;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [31:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [63:0] wire_16;
  assign wire_16 = L2End;
  wire [63:0] wire_17;
  wire [63:0] wire_18;
  wire [63:0] wire_18_0;
  wire [63:0] wire_18_1;
  assign wire_18 = wire_18_0|wire_18_1;
  wire [0:0] wire_19;
  wire [31:0] wire_20;
  wire [31:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [63:0] wire_24;
  assign wire_24 = L2Start;
  wire [0:0] wire_25;
  assign Output_1 = wire_25;
  wire [31:0] wire_26;
  wire [0:0] wire_27;
  wire [63:0] wire_28;
  assign wire_28 = L1Start;
  wire [31:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;

endmodule
