module _8bBitSelector (clk, rst, Number_1, Position, Number_2);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [63:0] Number_1;
  input  wire [7:0] Position;
  output  wire [63:0] Number_2;

  TC_Maker64 # (.UUID(64'd1312921996304714677 ^ UUID)) Maker64_0 (.in0(wire_11), .in1(wire_10), .in2(wire_6), .in3(wire_16), .in4(wire_19), .in5(wire_28), .in6(wire_34), .in7(wire_17), .out(wire_5));
  TC_Constant # (.UUID(64'd1341515457941498762 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_1 (.out(wire_25));
  TC_Constant # (.UUID(64'd4444718433828098485 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_2 (.out(wire_2));
  TC_Constant # (.UUID(64'd2003393661368942658 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_3 (.out(wire_23));
  TC_Constant # (.UUID(64'd3455227506599156849 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_4 (.out(wire_39));
  TC_Constant # (.UUID(64'd1052591411921414967 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_5 (.out(wire_29));
  TC_Constant # (.UUID(64'd205642527582532336 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5)) Constant8_6 (.out(wire_27));
  TC_Constant # (.UUID(64'd1274514892294560642 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h8)) Constant8_7 (.out(wire_15));
  TC_Constant # (.UUID(64'd668624861615954031 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_8 (.out(wire_36));
  TC_Splitter64 # (.UUID(64'd2747749493427573637 ^ UUID)) Splitter64_9 (.in(wire_35), .out0(wire_9), .out1(wire_8), .out2(wire_40), .out3(wire_3), .out4(wire_4), .out5(wire_38), .out6(wire_26), .out7(wire_1));
  TC_Maker32 # (.UUID(64'd1682693777870291492 ^ UUID)) Maker32_10 (.in0(wire_4), .in1(wire_38), .in2(wire_26), .in3(wire_1), .out(wire_32));
  TC_Splitter32 # (.UUID(64'd3460377708575970103 ^ UUID)) Splitter32_11 (.in(wire_32), .out0(wire_21), .out1(wire_30), .out2(wire_20), .out3(wire_41));
  TC_Maker16 # (.UUID(64'd139261840522345239 ^ UUID)) Maker16_12 (.in0(wire_40), .in1(wire_3), .out(wire_14));
  TC_Splitter16 # (.UUID(64'd4459133945486831877 ^ UUID)) Splitter16_13 (.in(wire_14), .out0(wire_18), .out1(wire_0));
  BitSelector # (.UUID(64'd813950653450767969 ^ UUID)) BitSelector_14 (.clk(clk), .rst(rst), .\8b_limit (wire_31), .\8b_Location (wire_25), .Number_1(wire_9), .Output(), .Number_2(wire_11));
  BitSelector # (.UUID(64'd2454877951581033315 ^ UUID)) BitSelector_15 (.clk(clk), .rst(rst), .\8b_limit (wire_22), .\8b_Location (wire_2), .Number_1(wire_8), .Output(wire_31), .Number_2(wire_10));
  BitSelector # (.UUID(64'd1509171945253359648 ^ UUID)) BitSelector_16 (.clk(clk), .rst(rst), .\8b_limit (wire_13), .\8b_Location (wire_23), .Number_1(wire_18), .Output(wire_22), .Number_2(wire_6));
  BitSelector # (.UUID(64'd4234163479417101366 ^ UUID)) BitSelector_17 (.clk(clk), .rst(rst), .\8b_limit (wire_12), .\8b_Location (wire_36), .Number_1(wire_0), .Output(wire_13), .Number_2(wire_16));
  BitSelector # (.UUID(64'd283819458352222539 ^ UUID)) BitSelector_18 (.clk(clk), .rst(rst), .\8b_limit (wire_37), .\8b_Location (wire_27), .Number_1(wire_21), .Output(wire_12), .Number_2(wire_19));
  BitSelector # (.UUID(64'd2850468475187288322 ^ UUID)) BitSelector_19 (.clk(clk), .rst(rst), .\8b_limit (wire_24), .\8b_Location (wire_29), .Number_1(wire_30), .Output(wire_37), .Number_2(wire_28));
  BitSelector # (.UUID(64'd3495643157198531230 ^ UUID)) BitSelector_20 (.clk(clk), .rst(rst), .\8b_limit (wire_33), .\8b_Location (wire_39), .Number_1(wire_20), .Output(wire_24), .Number_2(wire_34));
  BitSelector # (.UUID(64'd2860134298936815438 ^ UUID)) BitSelector_21 (.clk(clk), .rst(rst), .\8b_limit (wire_7), .\8b_Location (wire_15), .Number_1(wire_41), .Output(wire_33), .Number_2(wire_17));

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_3;
  wire [7:0] wire_4;
  wire [63:0] wire_5;
  assign Number_2 = wire_5;
  wire [7:0] wire_6;
  wire [7:0] wire_7;
  assign wire_7 = Position;
  wire [7:0] wire_8;
  wire [7:0] wire_9;
  wire [7:0] wire_10;
  wire [7:0] wire_11;
  wire [7:0] wire_12;
  wire [7:0] wire_13;
  wire [15:0] wire_14;
  wire [7:0] wire_15;
  wire [7:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_18;
  wire [7:0] wire_19;
  wire [7:0] wire_20;
  wire [7:0] wire_21;
  wire [7:0] wire_22;
  wire [7:0] wire_23;
  wire [7:0] wire_24;
  wire [7:0] wire_25;
  wire [7:0] wire_26;
  wire [7:0] wire_27;
  wire [7:0] wire_28;
  wire [7:0] wire_29;
  wire [7:0] wire_30;
  wire [7:0] wire_31;
  wire [31:0] wire_32;
  wire [7:0] wire_33;
  wire [7:0] wire_34;
  wire [63:0] wire_35;
  assign wire_35 = Number_1;
  wire [7:0] wire_36;
  wire [7:0] wire_37;
  wire [7:0] wire_38;
  wire [7:0] wire_39;
  wire [7:0] wire_40;
  wire [7:0] wire_41;

endmodule
