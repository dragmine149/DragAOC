module Day4Part1 (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_FileLoader # (.UUID(64'd1300333077211007914 ^ UUID), .DEFAULT_FILE_NAME("day4")) FileLoader_0 (.clk(clk), .rst(rst), .en(wire_57), .address({{56{1'b0}}, wire_65 }), .out(wire_14));
  TC_Constant # (.UUID(64'd614705877810942359 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_1 (.out(wire_57));
  TC_IndexerByte # (.UUID(64'd3259875342327518678 ^ UUID), .INDEX(64'd0)) IndexerByte_2 (.in(wire_14), .out(wire_7));
  TC_Constant # (.UUID(64'd2881157116684703501 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_3 (.out(wire_8));
  TC_IndexerByte # (.UUID(64'd3282167999629572026 ^ UUID), .INDEX(64'd0)) IndexerByte_4 (.in(wire_23), .out(wire_46));
  TC_IndexerByte # (.UUID(64'd344938491191684993 ^ UUID), .INDEX(64'd1)) IndexerByte_5 (.in(wire_23), .out(wire_64));
  TC_IndexerByte # (.UUID(64'd3057145202194435591 ^ UUID), .INDEX(64'd2)) IndexerByte_6 (.in(wire_23), .out(wire_33));
  TC_IndexerByte # (.UUID(64'd196694779505405906 ^ UUID), .INDEX(64'd3)) IndexerByte_7 (.in(wire_23), .out(wire_13));
  TC_IndexerByte # (.UUID(64'd195480252778983173 ^ UUID), .INDEX(64'd4)) IndexerByte_8 (.in(wire_23), .out(wire_58));
  TC_IndexerByte # (.UUID(64'd2249681588834216334 ^ UUID), .INDEX(64'd5)) IndexerByte_9 (.in(wire_23), .out(wire_39));
  TC_Maker64 # (.UUID(64'd2041678736802242094 ^ UUID)) Maker64_10 (.in0(wire_66), .in1(wire_67), .in2(wire_60), .in3(wire_45), .in4(wire_28), .in5(wire_61), .in6(8'd0), .in7(8'd0), .out(wire_23));
  TC_DelayLine # (.UUID(64'd1478884666127726678 ^ UUID), .BIT_WIDTH(64'd8)) DelayLine8_11 (.clk(clk), .rst(rst), .in(wire_40), .out(wire_65));
  TC_Constant # (.UUID(64'd4230246302748610089 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_12 (.out(wire_40));
  TC_IndexerByte # (.UUID(64'd3885874403913997322 ^ UUID), .INDEX(64'd1)) IndexerByte_13 (.in(wire_14), .out(wire_53));
  TC_IndexerByte # (.UUID(64'd2749811280805536878 ^ UUID), .INDEX(64'd2)) IndexerByte_14 (.in(wire_14), .out(wire_27));
  TC_IndexerByte # (.UUID(64'd3113000412030619556 ^ UUID), .INDEX(64'd3)) IndexerByte_15 (.in(wire_14), .out(wire_52));
  TC_IndexerByte # (.UUID(64'd3058128748266773168 ^ UUID), .INDEX(64'd4)) IndexerByte_16 (.in(wire_14), .out(wire_43));
  TC_IndexerByte # (.UUID(64'd3726479596336349432 ^ UUID), .INDEX(64'd5)) IndexerByte_17 (.in(wire_14), .out(wire_38));
  TC_Splitter64 # (.UUID(64'd1715894660434795144 ^ UUID)) Splitter64_18 (.in(wire_17), .out0(wire_25), .out1(wire_24), .out2(wire_0), .out3(wire_36), .out4(wire_26), .out5(wire_42), .out6(), .out7());
  TC_Switch # (.UUID(64'd3083524623901623221 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_19 (.en(wire_31), .in(wire_23), .out(wire_17));
  TC_Not # (.UUID(64'd1741588675539327596 ^ UUID), .BIT_WIDTH(64'd1)) Not_20 (.in(wire_4), .out(wire_31));
  TC_Counter # (.UUID(64'd2796646339049657840 ^ UUID), .BIT_WIDTH(64'd16), .count(16'd1)) Counter16_21 (.clk(clk), .rst(rst), .save(wire_56), .in(wire_6), .out(wire_6));
  TC_Not # (.UUID(64'd262671911581901502 ^ UUID), .BIT_WIDTH(64'd1)) Not_22 (.in(wire_62), .out(wire_56));
  TC_Halt # (.UUID(64'd2373505150995397943 ^ UUID), .HALT_MESSAGE("Upper limit reached")) Halt_23 (.clk(clk), .rst(rst), .en(wire_37));
  TC_Switch # (.UUID(64'd4386075278005230458 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_24 (.en(wire_31), .in(wire_5), .out(wire_37));
  TC_LessI # (.UUID(64'd3292654551045928704 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_25 (.in0(wire_1), .in1(wire_3), .out(wire_49));
  TC_LessI # (.UUID(64'd3747362352843898306 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_26 (.in0(wire_2), .in1(wire_1), .out(wire_12));
  TC_LessI # (.UUID(64'd4227878923150009143 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_27 (.in0(wire_16), .in1(wire_2), .out(wire_41));
  TC_LessI # (.UUID(64'd4090912352078921077 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_28 (.in0(wire_15), .in1(wire_16), .out(wire_18));
  TC_LessI # (.UUID(64'd2040532423834977934 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_29 (.in0(wire_20), .in1(wire_15), .out(wire_35));
  TC_Not # (.UUID(64'd366707461536672635 ^ UUID), .BIT_WIDTH(64'd1)) Not_30 (.in(wire_35), .out(wire_19));
  TC_Not # (.UUID(64'd2939040142042526066 ^ UUID), .BIT_WIDTH(64'd1)) Not_31 (.in(wire_18), .out(wire_34));
  TC_Not # (.UUID(64'd1398917821098271411 ^ UUID), .BIT_WIDTH(64'd1)) Not_32 (.in(wire_41), .out(wire_32));
  TC_Not # (.UUID(64'd3712273125459795596 ^ UUID), .BIT_WIDTH(64'd1)) Not_33 (.in(wire_12), .out(wire_54));
  TC_Not # (.UUID(64'd349618724439403530 ^ UUID), .BIT_WIDTH(64'd1)) Not_34 (.in(wire_49), .out(wire_68));
  TC_And # (.UUID(64'd949179814438959664 ^ UUID), .BIT_WIDTH(64'd1)) And_35 (.in0(wire_10), .in1(wire_11), .out(wire_47));
  TC_Switch # (.UUID(64'd3806424035603758608 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_36 (.en(wire_31), .in(wire_47), .out(wire_62));
  NotTick # (.UUID(64'd988254291887862844 ^ UUID)) NotTick_37 (.clk(clk), .rst(rst), .Output(wire_4));
  Cellz_2 # (.UUID(64'd2862707243587997049 ^ UUID)) Cellz_2_38 (.clk(clk), .rst(rst), .Increment(1'd0), .Overwrite(8'd0), .Global_Overwrite(1'd0), .Previous(8'd0), .Output(), .Increment_Next());
  Cellz_2 # (.UUID(64'd4552145864438261074 ^ UUID)) Cellz_2_39 (.clk(clk), .rst(rst), .Increment(1'd0), .Overwrite(8'd0), .Global_Overwrite(1'd0), .Previous(8'd0), .Output(), .Increment_Next());
  Cellz_2 # (.UUID(64'd3473631956184284865 ^ UUID)) Cellz_2_40 (.clk(clk), .rst(rst), .Increment(1'd0), .Overwrite(8'd0), .Global_Overwrite(1'd0), .Previous(8'd0), .Output(), .Increment_Next());
  Cellz_2 # (.UUID(64'd3264979902125614313 ^ UUID)) Cellz_2_41 (.clk(clk), .rst(rst), .Increment(1'd0), .Overwrite(8'd0), .Global_Overwrite(1'd0), .Previous(8'd0), .Output(), .Increment_Next());
  Cellz_2 # (.UUID(64'd848292611789013369 ^ UUID)) Cellz_2_42 (.clk(clk), .rst(rst), .Increment(1'd0), .Overwrite(8'd0), .Global_Overwrite(1'd0), .Previous(8'd0), .Output(), .Increment_Next());
  Cellz_2 # (.UUID(64'd4604342630189829407 ^ UUID)) Cellz_2_43 (.clk(clk), .rst(rst), .Increment(1'd0), .Overwrite(8'd0), .Global_Overwrite(1'd0), .Previous(8'd0), .Output(), .Increment_Next());
  ByteToNumber # (.UUID(64'd2290549341218488923 ^ UUID)) ByteToNumber_44 (.clk(clk), .rst(rst), .Input(wire_7), .Output(wire_66));
  ByteToNumber # (.UUID(64'd4267877789773175085 ^ UUID)) ByteToNumber_45 (.clk(clk), .rst(rst), .Input(wire_53), .Output(wire_67));
  ByteToNumber # (.UUID(64'd803095588841364073 ^ UUID)) ByteToNumber_46 (.clk(clk), .rst(rst), .Input(wire_27), .Output(wire_60));
  ByteToNumber # (.UUID(64'd677672594194363867 ^ UUID)) ByteToNumber_47 (.clk(clk), .rst(rst), .Input(wire_52), .Output(wire_45));
  ByteToNumber # (.UUID(64'd2617233141476735101 ^ UUID)) ByteToNumber_48 (.clk(clk), .rst(rst), .Input(wire_43), .Output(wire_28));
  ByteToNumber # (.UUID(64'd3235338507986847377 ^ UUID)) ByteToNumber_49 (.clk(clk), .rst(rst), .Input(wire_38), .Output(wire_61));
  _4beq # (.UUID(64'd4084947534873581742 ^ UUID)) _4beq_50 (.clk(clk), .rst(rst), .Input_1(wire_3), .Input_2(wire_1), .Output(wire_48));
  _4beq # (.UUID(64'd837930388802506938 ^ UUID)) _4beq_51 (.clk(clk), .rst(rst), .Input_1(wire_1), .Input_2(wire_2), .Output(wire_9));
  _4beq # (.UUID(64'd1001160964423906324 ^ UUID)) _4beq_52 (.clk(clk), .rst(rst), .Input_1(wire_2), .Input_2(wire_16), .Output(wire_59));
  _4beq # (.UUID(64'd4024915304172217312 ^ UUID)) _4beq_53 (.clk(clk), .rst(rst), .Input_1(wire_16), .Input_2(wire_15), .Output(wire_22));
  _4beq # (.UUID(64'd3801586074555563384 ^ UUID)) _4beq_54 (.clk(clk), .rst(rst), .Input_1(wire_15), .Input_2(wire_20), .Output(wire_55));
  OnOrOff # (.UUID(64'd2794213930716429597 ^ UUID)) OnOrOff_55 (.clk(clk), .rst(rst), .Input(wire_9), .Output(wire_10_3));
  OnOrOff # (.UUID(64'd321309780266364927 ^ UUID)) OnOrOff_56 (.clk(clk), .rst(rst), .Input(wire_59), .Output(wire_10_2));
  OnOrOff # (.UUID(64'd2791637861636592922 ^ UUID)) OnOrOff_57 (.clk(clk), .rst(rst), .Input(wire_22), .Output(wire_10_1));
  OnOrOff # (.UUID(64'd4363176194552780331 ^ UUID)) OnOrOff_58 (.clk(clk), .rst(rst), .Input(wire_55), .Output(wire_10_0));
  OnOrOff # (.UUID(64'd2565202741671842960 ^ UUID)) OnOrOff_59 (.clk(clk), .rst(rst), .Input(wire_48), .Output(wire_10_4));
  mand # (.UUID(64'd2743742951316189243 ^ UUID)) mand_60 (.clk(clk), .rst(rst), .Input_1(wire_68), .Input_2(wire_54), .Output(wire_29));
  mand # (.UUID(64'd2942067753606735184 ^ UUID)) mand_61 (.clk(clk), .rst(rst), .Input_1(wire_32), .Input_2(wire_34), .Output(wire_69));
  mand # (.UUID(64'd18958839450887314 ^ UUID)) mand_62 (.clk(clk), .rst(rst), .Input_1(wire_29), .Input_2(wire_63), .Output(wire_11));
  mand # (.UUID(64'd3212422335951933954 ^ UUID)) mand_63 (.clk(clk), .rst(rst), .Input_1(wire_69), .Input_2(wire_19), .Output(wire_63));
  RangeChecker # (.UUID(64'd2690237951565181585 ^ UUID)) RangeChecker_64 (.clk(clk), .rst(rst), .Input_1(wire_24), .Input_2(wire_1), .Input_3(wire_25), .Input_4(wire_3), .Input_5(wire_42), .Input_6(wire_20), .Input_7(wire_26), .Input_8(wire_15), .Input_9(wire_36), .Input_10(wire_16), .Input_11(wire_0), .Input_12(wire_2), .Output(wire_5));
  Cellz_2z_Dumb # (.UUID(64'd2574331762437855910 ^ UUID)) Cellz_2z_Dumb_65 (.clk(clk), .rst(rst), .Increment(1'd0), .Overwrite(8'd0), .Global_Overwrite(1'd0), .Output(), .Increment_Next());
  Cellz_2z_Dumb # (.UUID(64'd4175423220195224717 ^ UUID)) Cellz_2z_Dumb_66 (.clk(clk), .rst(rst), .Increment(wire_8), .Overwrite(wire_39), .Global_Overwrite(wire_4), .Output(wire_20), .Increment_Next(wire_50));
  Cellz_2z_Dumb # (.UUID(64'd356436453544593384 ^ UUID)) Cellz_2z_Dumb_67 (.clk(clk), .rst(rst), .Increment(wire_50), .Overwrite(wire_58), .Global_Overwrite(wire_4), .Output(wire_15), .Increment_Next(wire_51));
  Cellz_2z_Dumb # (.UUID(64'd2258755198707606320 ^ UUID)) Cellz_2z_Dumb_68 (.clk(clk), .rst(rst), .Increment(wire_51), .Overwrite(wire_13), .Global_Overwrite(wire_4), .Output(wire_16), .Increment_Next(wire_44));
  Cellz_2z_Dumb # (.UUID(64'd2804426362788026956 ^ UUID)) Cellz_2z_Dumb_69 (.clk(clk), .rst(rst), .Increment(wire_44), .Overwrite(wire_33), .Global_Overwrite(wire_4), .Output(wire_2), .Increment_Next(wire_21));
  Cellz_2z_Dumb # (.UUID(64'd381255555799844068 ^ UUID)) Cellz_2z_Dumb_70 (.clk(clk), .rst(rst), .Increment(wire_21), .Overwrite(wire_64), .Global_Overwrite(wire_4), .Output(wire_1), .Increment_Next(wire_30));
  Cellz_2z_Dumb # (.UUID(64'd2122555317477608146 ^ UUID)) Cellz_2z_Dumb_71 (.clk(clk), .rst(rst), .Increment(wire_30), .Overwrite(wire_46), .Global_Overwrite(wire_4), .Output(wire_3), .Increment_Next());

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [15:0] wire_6;
  wire [7:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_10_0;
  wire [0:0] wire_10_1;
  wire [0:0] wire_10_2;
  wire [0:0] wire_10_3;
  wire [0:0] wire_10_4;
  assign wire_10 = wire_10_0|wire_10_1|wire_10_2|wire_10_3|wire_10_4;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [7:0] wire_13;
  wire [63:0] wire_14;
  wire [7:0] wire_15;
  wire [7:0] wire_16;
  wire [63:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [7:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [63:0] wire_23;
  wire [7:0] wire_24;
  wire [7:0] wire_25;
  wire [7:0] wire_26;
  wire [7:0] wire_27;
  wire [7:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [7:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [7:0] wire_36;
  wire [0:0] wire_37;
  wire [7:0] wire_38;
  wire [7:0] wire_39;
  wire [7:0] wire_40;
  wire [0:0] wire_41;
  wire [7:0] wire_42;
  wire [7:0] wire_43;
  wire [0:0] wire_44;
  wire [7:0] wire_45;
  wire [7:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [7:0] wire_52;
  wire [7:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [7:0] wire_58;
  wire [0:0] wire_59;
  wire [7:0] wire_60;
  wire [7:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [7:0] wire_64;
  wire [7:0] wire_65;
  wire [7:0] wire_66;
  wire [7:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;

endmodule
