module Day4Part2 (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_FileLoader # (.UUID(64'd1300333077211007914 ^ UUID), .DEFAULT_FILE_NAME("day4")) FileLoader_0 (.clk(clk), .rst(rst), .en(wire_88), .address({{56{1'b0}}, wire_77 }), .out(wire_48));
  TC_Constant # (.UUID(64'd614705877810942359 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_1 (.out(wire_88));
  TC_IndexerByte # (.UUID(64'd3259875342327518678 ^ UUID), .INDEX(64'd0)) IndexerByte_2 (.in(wire_48), .out(wire_12));
  TC_Constant # (.UUID(64'd2881157116684703501 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_3 (.out(wire_50));
  TC_IndexerByte # (.UUID(64'd3282167999629572026 ^ UUID), .INDEX(64'd0)) IndexerByte_4 (.in(wire_41), .out(wire_82));
  TC_IndexerByte # (.UUID(64'd344938491191684993 ^ UUID), .INDEX(64'd1)) IndexerByte_5 (.in(wire_41), .out(wire_64));
  TC_IndexerByte # (.UUID(64'd3057145202194435591 ^ UUID), .INDEX(64'd2)) IndexerByte_6 (.in(wire_41), .out(wire_35));
  TC_IndexerByte # (.UUID(64'd196694779505405906 ^ UUID), .INDEX(64'd3)) IndexerByte_7 (.in(wire_41), .out(wire_40));
  TC_IndexerByte # (.UUID(64'd195480252778983173 ^ UUID), .INDEX(64'd4)) IndexerByte_8 (.in(wire_41), .out(wire_70));
  TC_IndexerByte # (.UUID(64'd2249681588834216334 ^ UUID), .INDEX(64'd5)) IndexerByte_9 (.in(wire_41), .out(wire_38));
  TC_Maker64 # (.UUID(64'd2041678736802242094 ^ UUID)) Maker64_10 (.in0(wire_46), .in1(wire_63), .in2(wire_79), .in3(wire_73), .in4(wire_55), .in5(wire_49), .in6(8'd0), .in7(8'd0), .out(wire_41));
  TC_DelayLine # (.UUID(64'd1478884666127726678 ^ UUID), .BIT_WIDTH(64'd8)) DelayLine8_11 (.clk(clk), .rst(rst), .in(wire_45), .out(wire_77));
  TC_Constant # (.UUID(64'd4230246302748610089 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_12 (.out(wire_45));
  TC_IndexerByte # (.UUID(64'd3885874403913997322 ^ UUID), .INDEX(64'd1)) IndexerByte_13 (.in(wire_48), .out(wire_57));
  TC_IndexerByte # (.UUID(64'd2749811280805536878 ^ UUID), .INDEX(64'd2)) IndexerByte_14 (.in(wire_48), .out(wire_58));
  TC_IndexerByte # (.UUID(64'd3113000412030619556 ^ UUID), .INDEX(64'd3)) IndexerByte_15 (.in(wire_48), .out(wire_52));
  TC_IndexerByte # (.UUID(64'd3058128748266773168 ^ UUID), .INDEX(64'd4)) IndexerByte_16 (.in(wire_48), .out(wire_29));
  TC_IndexerByte # (.UUID(64'd3726479596336349432 ^ UUID), .INDEX(64'd5)) IndexerByte_17 (.in(wire_48), .out(wire_84));
  TC_Splitter64 # (.UUID(64'd1715894660434795144 ^ UUID)) Splitter64_18 (.in(wire_65), .out0(wire_18), .out1(wire_56), .out2(wire_78), .out3(wire_67), .out4(wire_24), .out5(wire_33), .out6(), .out7());
  TC_Switch # (.UUID(64'd3083524623901623221 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_19 (.en(wire_15), .in(wire_41), .out(wire_65));
  TC_Not # (.UUID(64'd1741588675539327596 ^ UUID), .BIT_WIDTH(64'd1)) Not_20 (.in(wire_14), .out(wire_15));
  TC_Counter # (.UUID(64'd2796646339049657840 ^ UUID), .BIT_WIDTH(64'd16), .count(16'd1)) Counter16_21 (.clk(clk), .rst(rst), .save(wire_71), .in(wire_23), .out(wire_23));
  TC_Not # (.UUID(64'd262671911581901502 ^ UUID), .BIT_WIDTH(64'd1)) Not_22 (.in(wire_86), .out(wire_71));
  TC_Halt # (.UUID(64'd2373505150995397943 ^ UUID), .HALT_MESSAGE("Upper limit reached")) Halt_23 (.clk(clk), .rst(rst), .en(wire_16));
  TC_Switch # (.UUID(64'd4386075278005230458 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_24 (.en(wire_15), .in(wire_81), .out(wire_16));
  TC_LessI # (.UUID(64'd3292654551045928704 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_25 (.in0(wire_3), .in1(wire_30), .out(wire_68));
  TC_LessI # (.UUID(64'd3747362352843898306 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_26 (.in0(wire_9), .in1(wire_3), .out(wire_53));
  TC_LessI # (.UUID(64'd4227878923150009143 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_27 (.in0(wire_13), .in1(wire_9), .out(wire_62));
  TC_LessI # (.UUID(64'd4090912352078921077 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_28 (.in0(wire_11), .in1(wire_13), .out(wire_66));
  TC_LessI # (.UUID(64'd2040532423834977934 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_29 (.in0(wire_28), .in1(wire_11), .out(wire_60));
  TC_Not # (.UUID(64'd366707461536672635 ^ UUID), .BIT_WIDTH(64'd1)) Not_30 (.in(wire_60), .out(wire_32));
  TC_Not # (.UUID(64'd2939040142042526066 ^ UUID), .BIT_WIDTH(64'd1)) Not_31 (.in(wire_66), .out(wire_43));
  TC_Not # (.UUID(64'd1398917821098271411 ^ UUID), .BIT_WIDTH(64'd1)) Not_32 (.in(wire_62), .out(wire_83));
  TC_Not # (.UUID(64'd3712273125459795596 ^ UUID), .BIT_WIDTH(64'd1)) Not_33 (.in(wire_53), .out(wire_47));
  TC_Not # (.UUID(64'd349618724439403530 ^ UUID), .BIT_WIDTH(64'd1)) Not_34 (.in(wire_68), .out(wire_54));
  TC_And # (.UUID(64'd949179814438959664 ^ UUID), .BIT_WIDTH(64'd1)) And_35 (.in0(wire_4), .in1(wire_75), .out(wire_39));
  TC_Switch # (.UUID(64'd3806424035603758608 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_36 (.en(wire_15), .in(wire_39), .out(wire_86));
  TC_Switch # (.UUID(64'd3815757842053566393 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_37 (.en(wire_89), .in(wire_50), .out(wire_72));
  TC_Not # (.UUID(64'd4517909894909000332 ^ UUID), .BIT_WIDTH(64'd1)) Not_38 (.in(wire_85), .out(wire_89));
  TC_DelayLine # (.UUID(64'd1998668017909422993 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_39 (.clk(clk), .rst(rst), .in(wire_26), .out(wire_85));
  TC_DelayLine # (.UUID(64'd2142609526691430932 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_40 (.clk(clk), .rst(rst), .in(wire_44), .out(wire_87));
  NotTick # (.UUID(64'd988254291887862844 ^ UUID)) NotTick_41 (.clk(clk), .rst(rst), .Output(wire_14));
  ByteToNumber # (.UUID(64'd2290549341218488923 ^ UUID)) ByteToNumber_42 (.clk(clk), .rst(rst), .Input(wire_12), .Output(wire_46));
  ByteToNumber # (.UUID(64'd4267877789773175085 ^ UUID)) ByteToNumber_43 (.clk(clk), .rst(rst), .Input(wire_57), .Output(wire_63));
  ByteToNumber # (.UUID(64'd803095588841364073 ^ UUID)) ByteToNumber_44 (.clk(clk), .rst(rst), .Input(wire_58), .Output(wire_79));
  ByteToNumber # (.UUID(64'd677672594194363867 ^ UUID)) ByteToNumber_45 (.clk(clk), .rst(rst), .Input(wire_52), .Output(wire_73));
  ByteToNumber # (.UUID(64'd2617233141476735101 ^ UUID)) ByteToNumber_46 (.clk(clk), .rst(rst), .Input(wire_29), .Output(wire_55));
  ByteToNumber # (.UUID(64'd3235338507986847377 ^ UUID)) ByteToNumber_47 (.clk(clk), .rst(rst), .Input(wire_84), .Output(wire_49));
  mand # (.UUID(64'd2743742951316189243 ^ UUID)) mand_48 (.clk(clk), .rst(rst), .Input_1(wire_54), .Input_2(wire_47), .Output(wire_37));
  mand # (.UUID(64'd2942067753606735184 ^ UUID)) mand_49 (.clk(clk), .rst(rst), .Input_1(wire_83), .Input_2(wire_43), .Output(wire_34));
  mand # (.UUID(64'd18958839450887314 ^ UUID)) mand_50 (.clk(clk), .rst(rst), .Input_1(wire_37), .Input_2(wire_80), .Output(wire_75));
  mand # (.UUID(64'd3212422335951933954 ^ UUID)) mand_51 (.clk(clk), .rst(rst), .Input_1(wire_34), .Input_2(wire_32), .Output(wire_80));
  RangeChecker # (.UUID(64'd2690237951565181585 ^ UUID)) RangeChecker_52 (.clk(clk), .rst(rst), .Input_1(wire_56), .Input_2(wire_3), .Input_3(wire_18), .Input_4(wire_30), .Input_5(wire_33), .Input_6(wire_28), .Input_7(wire_24), .Input_8(wire_11), .Input_9(wire_67), .Input_10(wire_13), .Input_11(wire_78), .Input_12(wire_9), .Output(wire_81));
  Cellz_2 # (.UUID(64'd2681121728217391920 ^ UUID)) Cellz_2_53 (.clk(clk), .rst(rst), .Increment(wire_22), .Overwrite(wire_82), .Global_Overwrite(wire_14), .Previous(8'd0), .Output(wire_30), .Increment_Next());
  Cellz_2 # (.UUID(64'd3469695128675857344 ^ UUID)) Cellz_2_54 (.clk(clk), .rst(rst), .Increment(wire_27), .Overwrite(wire_64), .Global_Overwrite(wire_14), .Previous(wire_30), .Output(wire_3), .Increment_Next(wire_22));
  Cellz_2 # (.UUID(64'd2464365340593423882 ^ UUID)) Cellz_2_55 (.clk(clk), .rst(rst), .Increment(wire_61), .Overwrite(wire_35), .Global_Overwrite(wire_14), .Previous(wire_3), .Output(wire_9), .Increment_Next(wire_27));
  Cellz_2 # (.UUID(64'd403371948968645324 ^ UUID)) Cellz_2_56 (.clk(clk), .rst(rst), .Increment(wire_5), .Overwrite(wire_40), .Global_Overwrite(wire_14), .Previous(wire_9), .Output(wire_13), .Increment_Next(wire_61));
  Cellz_2 # (.UUID(64'd1534890721647203275 ^ UUID)) Cellz_2_57 (.clk(clk), .rst(rst), .Increment(wire_0), .Overwrite(wire_70), .Global_Overwrite(wire_14), .Previous(wire_13), .Output(wire_11), .Increment_Next(wire_5));
  Cellz_2 # (.UUID(64'd2165210612851354234 ^ UUID)) Cellz_2_58 (.clk(clk), .rst(rst), .Increment(wire_72), .Overwrite(wire_38), .Global_Overwrite(wire_14), .Previous(wire_11), .Output(wire_28), .Increment_Next(wire_0));
  OnOrOff # (.UUID(64'd129879025491825736 ^ UUID)) OnOrOff_59 (.clk(clk), .rst(rst), .Input(wire_22), .Output(wire_44_1));
  OnOrOff # (.UUID(64'd2069905977387596 ^ UUID)) OnOrOff_60 (.clk(clk), .rst(rst), .Input(wire_27), .Output(wire_44_0));
  OnOrOff # (.UUID(64'd4020034695276023527 ^ UUID)) OnOrOff_61 (.clk(clk), .rst(rst), .Input(wire_61), .Output(wire_26_2));
  OnOrOff # (.UUID(64'd3681849683264036923 ^ UUID)) OnOrOff_62 (.clk(clk), .rst(rst), .Input(wire_5), .Output(wire_26_1));
  OnOrOff # (.UUID(64'd1477728482954482203 ^ UUID)) OnOrOff_63 (.clk(clk), .rst(rst), .Input(wire_0), .Output(wire_26_0));
  OnOrOff # (.UUID(64'd2385286065099818749 ^ UUID)) OnOrOff_64 (.clk(clk), .rst(rst), .Input(wire_87), .Output(wire_26_3));
  _4beq # (.UUID(64'd2686310176453389258 ^ UUID)) _4beq_65 (.clk(clk), .rst(rst), .Input_1(wire_30), .Input_2(wire_3), .Output(wire_20));
  _4beq # (.UUID(64'd3482198435573910046 ^ UUID)) _4beq_66 (.clk(clk), .rst(rst), .Input_1(wire_3), .Input_2(wire_9), .Output(wire_25));
  _4beq # (.UUID(64'd3633788093279011507 ^ UUID)) _4beq_67 (.clk(clk), .rst(rst), .Input_1(wire_9), .Input_2(wire_13), .Output(wire_6));
  _4beq # (.UUID(64'd628268869804084334 ^ UUID)) _4beq_68 (.clk(clk), .rst(rst), .Input_1(wire_13), .Input_2(wire_11), .Output(wire_2));
  _4beq # (.UUID(64'd258847199856683304 ^ UUID)) _4beq_69 (.clk(clk), .rst(rst), .Input_1(wire_11), .Input_2(wire_28), .Output(wire_36));
  mand # (.UUID(64'd4560922881634669559 ^ UUID)) mand_70 (.clk(clk), .rst(rst), .Input_1(wire_20), .Input_2(wire_25), .Output(wire_17));
  TC_Not # (.UUID(64'd1902849945845820013 ^ UUID), .BIT_WIDTH(64'd1)) Not_71 (.in(wire_17), .out(wire_8));
  TC_Switch # (.UUID(64'd1974696222326850979 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_72 (.en(wire_8), .in(wire_20), .out(wire_10));
  OnOrOff # (.UUID(64'd2452945791868363870 ^ UUID)) OnOrOff_73 (.clk(clk), .rst(rst), .Input(wire_10), .Output(wire_4_2));
  mand # (.UUID(64'd3210724723724383364 ^ UUID)) mand_74 (.clk(clk), .rst(rst), .Input_1(wire_25), .Input_2(wire_6), .Output(wire_1));
  OnOrOff # (.UUID(64'd3988557037053602878 ^ UUID)) OnOrOff_75 (.clk(clk), .rst(rst), .Input(wire_21), .Output(wire_4_0));
  mand # (.UUID(64'd4238428015963384406 ^ UUID)) mand_76 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_2), .Output(wire_7));
  OnOrOff # (.UUID(64'd129812558163807238 ^ UUID)) OnOrOff_77 (.clk(clk), .rst(rst), .Input(wire_59), .Output(wire_4_1));
  mand # (.UUID(64'd3884660465656345454 ^ UUID)) mand_78 (.clk(clk), .rst(rst), .Input_1(wire_2), .Input_2(wire_36), .Output(wire_31));
  OnOrOff # (.UUID(64'd4219029386912714114 ^ UUID)) OnOrOff_79 (.clk(clk), .rst(rst), .Input(wire_42), .Output(wire_4_3));
  TC_Not # (.UUID(64'd4407995118227157989 ^ UUID), .BIT_WIDTH(64'd1)) Not_80 (.in(wire_31), .out(wire_51));
  TC_Switch # (.UUID(64'd1043627780545808567 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_81 (.en(wire_51), .in(wire_36), .out(wire_74));
  OnOrOff # (.UUID(64'd3015556203815749349 ^ UUID)) OnOrOff_82 (.clk(clk), .rst(rst), .Input(wire_74), .Output(wire_4_4));
  mand # (.UUID(64'd2496340798535357342 ^ UUID)) mand_83 (.clk(clk), .rst(rst), .Input_1(wire_69), .Input_2(wire_2), .Output(wire_42));
  mand # (.UUID(64'd108201680620660856 ^ UUID)) mand_84 (.clk(clk), .rst(rst), .Input_1(wire_76), .Input_2(wire_6), .Output(wire_59));
  mand # (.UUID(64'd299826000917452259 ^ UUID)) mand_85 (.clk(clk), .rst(rst), .Input_1(wire_19), .Input_2(wire_25), .Output(wire_21));
  mNOR # (.UUID(64'd2327488911447820817 ^ UUID)) mNOR_86 (.clk(clk), .rst(rst), .Input_1(wire_1), .Input_2(wire_17), .Output(wire_19));
  mNOR # (.UUID(64'd3660306186097943822 ^ UUID)) mNOR_87 (.clk(clk), .rst(rst), .Input_1(wire_7), .Input_2(wire_1), .Output(wire_76));
  mNOR # (.UUID(64'd3891289534251045762 ^ UUID)) mNOR_88 (.clk(clk), .rst(rst), .Input_1(wire_31), .Input_2(wire_7), .Output(wire_69));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [7:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_4_0;
  wire [0:0] wire_4_1;
  wire [0:0] wire_4_2;
  wire [0:0] wire_4_3;
  wire [0:0] wire_4_4;
  assign wire_4 = wire_4_0|wire_4_1|wire_4_2|wire_4_3|wire_4_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [7:0] wire_9;
  wire [0:0] wire_10;
  wire [7:0] wire_11;
  wire [7:0] wire_12;
  wire [7:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [7:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [15:0] wire_23;
  wire [7:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_26_0;
  wire [0:0] wire_26_1;
  wire [0:0] wire_26_2;
  wire [0:0] wire_26_3;
  assign wire_26 = wire_26_0|wire_26_1|wire_26_2|wire_26_3;
  wire [0:0] wire_27;
  wire [7:0] wire_28;
  wire [7:0] wire_29;
  wire [7:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [7:0] wire_33;
  wire [0:0] wire_34;
  wire [7:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [7:0] wire_38;
  wire [0:0] wire_39;
  wire [7:0] wire_40;
  wire [63:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_44_0;
  wire [0:0] wire_44_1;
  assign wire_44 = wire_44_0|wire_44_1;
  wire [7:0] wire_45;
  wire [7:0] wire_46;
  wire [0:0] wire_47;
  wire [63:0] wire_48;
  wire [7:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [7:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [7:0] wire_55;
  wire [7:0] wire_56;
  wire [7:0] wire_57;
  wire [7:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [7:0] wire_63;
  wire [7:0] wire_64;
  wire [63:0] wire_65;
  wire [0:0] wire_66;
  wire [7:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;
  wire [7:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [7:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [7:0] wire_77;
  wire [7:0] wire_78;
  wire [7:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [7:0] wire_82;
  wire [0:0] wire_83;
  wire [7:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;

endmodule
