module Day1Part1 (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_Register # (.UUID(64'd4178573859148191576 ^ UUID), .BIT_WIDTH(64'd64)) Register64_0 (.clk(clk), .rst(rst), .load(wire_37), .save(wire_28), .in(wire_24), .out(wire_23));
  TC_Add # (.UUID(64'd359763711881990385 ^ UUID), .BIT_WIDTH(64'd64)) Add64_1 (.in0({{56{1'b0}}, wire_29 }), .in1(wire_23), .ci(1'd0), .out(wire_24), .co());
  TC_Equal # (.UUID(64'd928735983604669128 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_2 (.in0(wire_29), .in1(wire_10), .out(wire_33));
  TC_Constant # (.UUID(64'd2218857169047162011 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h9)) Constant8_3 (.out(wire_10));
  TC_Counter # (.UUID(64'd1097574418592050277 ^ UUID), .BIT_WIDTH(64'd64), .count(64'd1)) Counter64_4 (.clk(clk), .rst(rst), .save(wire_5), .in(wire_30), .out(wire_30));
  TC_Register # (.UUID(64'd2413979704567083807 ^ UUID), .BIT_WIDTH(64'd64)) Register64_5 (.clk(clk), .rst(rst), .load(wire_15), .save(wire_26), .in(wire_21), .out(wire_4));
  TC_Constant # (.UUID(64'd2793433701128027946 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFFFFFFFFFFFFFFFF)) Constant64_6 (.out(wire_25));
  TC_Constant # (.UUID(64'd1184275376460161862 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_7 (.out(wire_15));
  TC_Not # (.UUID(64'd4603214268349776896 ^ UUID), .BIT_WIDTH(64'd1)) Not_8 (.in(wire_9), .out(wire_26));
  TC_Mux # (.UUID(64'd3836885967411031723 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_9 (.sel(wire_9), .in0(wire_25), .in1(wire_23), .out(wire_6));
  TC_DelayLine # (.UUID(64'd2178678318095205493 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_10 (.clk(clk), .rst(rst), .in(wire_36), .out(wire_19));
  TC_Not # (.UUID(64'd1630915932547760616 ^ UUID), .BIT_WIDTH(64'd1)) Not_11 (.in(wire_5), .out(wire_28));
  TC_Constant # (.UUID(64'd2213483610403812941 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_12 (.out(wire_37));
  TC_Not # (.UUID(64'd2394884979716713933 ^ UUID), .BIT_WIDTH(64'd1)) Not_13 (.in(wire_9), .out(wire_12));
  TC_Ram # (.UUID(64'd811351278422078506 ^ UUID), .WORD_WIDTH(64'd64), .WORD_COUNT(64'd1250)) Ram_14 (.clk(clk), .rst(rst), .load(wire_22), .save(wire_17), .address(wire_27[31:0]), .in0(wire_7), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_31), .out1(), .out2(), .out3());
  TC_FileLoader # (.UUID(64'd2193553924715941358 ^ UUID), .DEFAULT_FILE_NAME("day1")) FileLoader_15 (.clk(clk), .rst(rst), .en(wire_38), .address(wire_6), .out(wire_21));
  TC_Constant # (.UUID(64'd3595939561111802633 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_16 (.out(wire_38));
  TC_Switch # (.UUID(64'd3013778101405626680 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_17 (.en(wire_0), .in(wire_28), .out(wire_17));
  TC_Switch # (.UUID(64'd3957714978086000962 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_18 (.en(wire_0), .in(wire_30), .out(wire_27_1));
  TC_Switch # (.UUID(64'd4006497041254316547 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_19 (.en(wire_0), .in(wire_2), .out(wire_7));
  TC_LessU # (.UUID(64'd2412733997253528222 ^ UUID), .BIT_WIDTH(64'd64)) LessU64_20 (.in0(wire_23), .in1(wire_4), .out(wire_0));
  TC_Register # (.UUID(64'd1998148612828582261 ^ UUID), .BIT_WIDTH(64'd64)) Register64_21 (.clk(clk), .rst(rst), .load(wire_20), .save(wire_22), .in(wire_39), .out(wire_3));
  TC_Add # (.UUID(64'd3023020307212303517 ^ UUID), .BIT_WIDTH(64'd64)) Add64_22 (.in0(wire_8), .in1(wire_3), .ci(1'd0), .out(wire_39), .co());
  TC_Constant # (.UUID(64'd1388399570672712544 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_23 (.out(wire_20));
  TC_Counter # (.UUID(64'd1973994861164209717 ^ UUID), .BIT_WIDTH(64'd64), .count(64'd1)) Counter64_24 (.clk(clk), .rst(rst), .save(wire_18), .in(wire_16), .out(wire_16));
  TC_Not # (.UUID(64'd927835141595733835 ^ UUID), .BIT_WIDTH(64'd1)) Not_25 (.in(wire_0), .out(wire_35));
  TC_FileLoader # (.UUID(64'd1289831107320614410 ^ UUID), .DEFAULT_FILE_NAME("day1_test_1")) FileLoader_26 (.clk(clk), .rst(rst), .en(1'd0), .address(64'd0), .out());
  TC_Register # (.UUID(64'd2632168926008665082 ^ UUID), .BIT_WIDTH(64'd64)) Register64_27 (.clk(clk), .rst(rst), .load(wire_13), .save(wire_11), .in(wire_30), .out(wire_1));
  TC_Switch # (.UUID(64'd2600677178569538476 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_28 (.en(wire_34), .in(wire_35), .out(wire_11));
  TC_DelayLine # (.UUID(64'd3616072873250103679 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_29 (.clk(clk), .rst(rst), .in(wire_0), .out(wire_34));
  TC_Constant # (.UUID(64'd1666034379207229566 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_30 (.out(wire_13));
  TC_Not # (.UUID(64'd101522584180394033 ^ UUID), .BIT_WIDTH(64'd1)) Not_31 (.in(wire_22), .out(wire_18));
  TC_Equal # (.UUID(64'd4073392919419213019 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_32 (.in0(wire_16), .in1(wire_1), .out(wire_14));
  TC_Halt # (.UUID(64'd805079572016111755 ^ UUID), .HALT_MESSAGE("Program finished!")) Halt_33 (.clk(clk), .rst(rst), .en(wire_32));
  TC_Switch # (.UUID(64'd1270767012348834115 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_34 (.en(wire_22), .in(wire_14), .out(wire_32));
  BytesToNumbers # (.UUID(64'd4206582659042050133 ^ UUID)) BytesToNumbers_35 (.clk(clk), .rst(rst), .Carry(wire_19), .\Input_(64b) (wire_21), .Offset(wire_29), .\Output_(8b) (wire_2));
  _64zmany # (.UUID(64'd3133133748172620224 ^ UUID)) _64zmany_36 (.clk(clk), .rst(rst), .Input(wire_4), .Output(wire_9));
  flippedzm64bzmswitch # (.UUID(64'd1985891020947270661 ^ UUID)) flippedzm64bzmswitch_37 (.clk(clk), .rst(rst), .Input_1(wire_2), .Input_2(wire_33), .Output(wire_36));
  OnOrOff # (.UUID(64'd1600200685999643413 ^ UUID)) OnOrOff_38 (.clk(clk), .rst(rst), .Input(wire_33), .Output(wire_5_1));
  OnOrOff # (.UUID(64'd946715927199943045 ^ UUID)) OnOrOff_39 (.clk(clk), .rst(rst), .Input(wire_12), .Output(wire_5_0));
  Div3z_roundz_minusz_2 # (.UUID(64'd2501588780423282301 ^ UUID)) Div3z_roundz_minusz_2_40 (.clk(clk), .rst(rst), .Input(wire_31), .Output(wire_8));
  flippedzm64bzmswitch # (.UUID(64'd380343949002747622 ^ UUID)) flippedzm64bzmswitch_41 (.clk(clk), .rst(rst), .Input_1(wire_16), .Input_2(wire_35), .Output(wire_27_0));
  _64zmany # (.UUID(64'd2095873869615652318 ^ UUID)) _64zmany_42 (.clk(clk), .rst(rst), .Input(wire_1), .Output(wire_22));

  wire [0:0] wire_0;
  wire [63:0] wire_1;
  wire [63:0] wire_2;
  wire [63:0] wire_3;
  wire [63:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_5_0;
  wire [0:0] wire_5_1;
  assign wire_5 = wire_5_0|wire_5_1;
  wire [63:0] wire_6;
  wire [63:0] wire_7;
  wire [63:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [63:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [63:0] wire_19;
  wire [0:0] wire_20;
  wire [63:0] wire_21;
  wire [0:0] wire_22;
  wire [63:0] wire_23;
  wire [63:0] wire_24;
  wire [63:0] wire_25;
  wire [0:0] wire_26;
  wire [63:0] wire_27;
  wire [63:0] wire_27_0;
  wire [63:0] wire_27_1;
  assign wire_27 = wire_27_0|wire_27_1;
  wire [0:0] wire_28;
  wire [7:0] wire_29;
  wire [63:0] wire_30;
  wire [63:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [63:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [63:0] wire_39;

endmodule
