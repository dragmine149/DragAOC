module _8bNewLine (clk, rst, Input, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [63:0] Input;
  output  wire [7:0] Output;

  TC_Splitter64 # (.UUID(64'd3895924655864399812 ^ UUID)) Splitter64_0 (.in(wire_33), .out0(wire_16), .out1(wire_29), .out2(wire_0), .out3(wire_25), .out4(wire_14), .out5(wire_18), .out6(wire_7), .out7(wire_4));
  TC_Constant # (.UUID(64'd4508484919927074214 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_1 (.out(wire_48));
  TC_Constant # (.UUID(64'd2940396106940393774 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_2 (.out(wire_34));
  TC_Constant # (.UUID(64'd2157846558509232567 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_3 (.out(wire_27));
  TC_Constant # (.UUID(64'd205443766022644447 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_4 (.out(wire_37));
  TC_Constant # (.UUID(64'd3997912978879554374 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_5 (.out(wire_8));
  TC_Constant # (.UUID(64'd1105061765928732701 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5)) Constant8_6 (.out(wire_12));
  TC_Constant # (.UUID(64'd3801071687550733994 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_7 (.out(wire_39));
  TC_Constant # (.UUID(64'd1069872183118685998 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h8)) Constant8_8 (.out(wire_19));
  TC_Switch # (.UUID(64'd1747830201043249029 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_9 (.en(wire_44), .in(wire_6), .out(wire_35_0));
  TC_Not # (.UUID(64'd221836309478339864 ^ UUID), .BIT_WIDTH(64'd1)) Not_10 (.in(wire_11), .out(wire_44));
  newlineDetector # (.UUID(64'd1825159156690185713 ^ UUID)) newlineDetector_11 (.clk(clk), .rst(rst), .\Number_a._-45 (wire_25), .Index(wire_39), .Output(wire_5));
  newlineDetector # (.UUID(64'd3151820960339829815 ^ UUID)) newlineDetector_12 (.clk(clk), .rst(rst), .\Number_a._-45 (wire_0), .Index(wire_27), .Output(wire_38));
  newlineDetector # (.UUID(64'd2029869491286418204 ^ UUID)) newlineDetector_13 (.clk(clk), .rst(rst), .\Number_a._-45 (wire_29), .Index(wire_34), .Output(wire_13));
  newlineDetector # (.UUID(64'd3595269546581004239 ^ UUID)) newlineDetector_14 (.clk(clk), .rst(rst), .\Number_a._-45 (wire_16), .Index(wire_48), .Output(wire_2));
  newlineDetector # (.UUID(64'd1560030053312584685 ^ UUID)) newlineDetector_15 (.clk(clk), .rst(rst), .\Number_a._-45 (wire_7), .Index(wire_37), .Output(wire_28));
  newlineDetector # (.UUID(64'd3216684887509029446 ^ UUID)) newlineDetector_16 (.clk(clk), .rst(rst), .\Number_a._-45 (wire_18), .Index(wire_8), .Output(wire_3));
  newlineDetector # (.UUID(64'd4105934187413501361 ^ UUID)) newlineDetector_17 (.clk(clk), .rst(rst), .\Number_a._-45 (wire_14), .Index(wire_12), .Output(wire_1));
  newlineDetector # (.UUID(64'd2836405010755731853 ^ UUID)) newlineDetector_18 (.clk(clk), .rst(rst), .\Number_a._-45 (8'd0), .Index(8'd0), .Output(wire_41));
  _8zmany # (.UUID(64'd714338964245414581 ^ UUID)) _8zmany_19 (.clk(clk), .rst(rst), .Input(wire_2), .Output(wire_11));
  flippedzm8bzmswitch # (.UUID(64'd3830625961092996974 ^ UUID)) flippedzm8bzmswitch_20 (.clk(clk), .rst(rst), .Input_1(wire_2), .Input_2(wire_11), .Output(wire_35_1));
  TC_Not # (.UUID(64'd3002566734186577845 ^ UUID), .BIT_WIDTH(64'd1)) Not_21 (.in(wire_43), .out(wire_47));
  _8zmany # (.UUID(64'd1242029082602216693 ^ UUID)) _8zmany_22 (.clk(clk), .rst(rst), .Input(wire_13), .Output(wire_43));
  flippedzm8bzmswitch # (.UUID(64'd671695906598487034 ^ UUID)) flippedzm8bzmswitch_23 (.clk(clk), .rst(rst), .Input_1(wire_13), .Input_2(wire_43), .Output(wire_6_0));
  TC_Not # (.UUID(64'd1031601450290599409 ^ UUID), .BIT_WIDTH(64'd1)) Not_24 (.in(wire_17), .out(wire_46));
  _8zmany # (.UUID(64'd498655951945221264 ^ UUID)) _8zmany_25 (.clk(clk), .rst(rst), .Input(wire_38), .Output(wire_17));
  flippedzm8bzmswitch # (.UUID(64'd3406251113222130696 ^ UUID)) flippedzm8bzmswitch_26 (.clk(clk), .rst(rst), .Input_1(wire_38), .Input_2(wire_17), .Output(wire_36_0));
  TC_Not # (.UUID(64'd3679236801590722114 ^ UUID), .BIT_WIDTH(64'd1)) Not_27 (.in(wire_9), .out(wire_40));
  _8zmany # (.UUID(64'd3483365898671451887 ^ UUID)) _8zmany_28 (.clk(clk), .rst(rst), .Input(wire_5), .Output(wire_9));
  flippedzm8bzmswitch # (.UUID(64'd828850458229468365 ^ UUID)) flippedzm8bzmswitch_29 (.clk(clk), .rst(rst), .Input_1(wire_5), .Input_2(wire_9), .Output(wire_21_0));
  TC_Not # (.UUID(64'd2992545497868994766 ^ UUID), .BIT_WIDTH(64'd1)) Not_30 (.in(wire_32), .out(wire_23));
  _8zmany # (.UUID(64'd338285859100298700 ^ UUID)) _8zmany_31 (.clk(clk), .rst(rst), .Input(wire_1), .Output(wire_32));
  flippedzm8bzmswitch # (.UUID(64'd430241336298863432 ^ UUID)) flippedzm8bzmswitch_32 (.clk(clk), .rst(rst), .Input_1(wire_1), .Input_2(wire_32), .Output(wire_24_1));
  TC_Not # (.UUID(64'd2860553486456588788 ^ UUID), .BIT_WIDTH(64'd1)) Not_33 (.in(wire_26), .out(wire_15));
  _8zmany # (.UUID(64'd1750922629869402274 ^ UUID)) _8zmany_34 (.clk(clk), .rst(rst), .Input(wire_3), .Output(wire_26));
  flippedzm8bzmswitch # (.UUID(64'd261758794925260442 ^ UUID)) flippedzm8bzmswitch_35 (.clk(clk), .rst(rst), .Input_1(wire_3), .Input_2(wire_26), .Output(wire_22_0));
  TC_Not # (.UUID(64'd4590207191988151946 ^ UUID), .BIT_WIDTH(64'd1)) Not_36 (.in(wire_31), .out(wire_45));
  _8zmany # (.UUID(64'd1199315494658476821 ^ UUID)) _8zmany_37 (.clk(clk), .rst(rst), .Input(wire_28), .Output(wire_31));
  flippedzm8bzmswitch # (.UUID(64'd1457447456130014861 ^ UUID)) flippedzm8bzmswitch_38 (.clk(clk), .rst(rst), .Input_1(wire_28), .Input_2(wire_31), .Output(wire_10_1));
  TC_Not # (.UUID(64'd4476199958934872118 ^ UUID), .BIT_WIDTH(64'd1)) Not_39 (.in(wire_42), .out(wire_20));
  _8zmany # (.UUID(64'd2982169432180539901 ^ UUID)) _8zmany_40 (.clk(clk), .rst(rst), .Input(wire_41), .Output(wire_42));
  flippedzm8bzmswitch # (.UUID(64'd1986627394009335625 ^ UUID)) flippedzm8bzmswitch_41 (.clk(clk), .rst(rst), .Input_1(wire_41), .Input_2(wire_42), .Output(wire_30_1));
  TC_Switch # (.UUID(64'd2603706298106505537 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_42 (.en(wire_47), .in(wire_36), .out(wire_6_1));
  TC_Switch # (.UUID(64'd3135166035656658902 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_43 (.en(wire_46), .in(wire_21), .out(wire_36_1));
  TC_Switch # (.UUID(64'd3649895533361336479 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_44 (.en(wire_40), .in(wire_24), .out(wire_21_1));
  TC_Switch # (.UUID(64'd350126338011032993 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_45 (.en(wire_23), .in(wire_22), .out(wire_24_0));
  TC_Switch # (.UUID(64'd348013912476434600 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_46 (.en(wire_15), .in(wire_10), .out(wire_22_1));
  TC_Switch # (.UUID(64'd3605896724580726997 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_47 (.en(wire_45), .in(wire_30), .out(wire_10_0));
  TC_Switch # (.UUID(64'd1763960916745122359 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_48 (.en(wire_20), .in(wire_19), .out(wire_30_0));

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_3;
  wire [7:0] wire_4;
  wire [7:0] wire_5;
  wire [7:0] wire_6;
  wire [7:0] wire_6_0;
  wire [7:0] wire_6_1;
  assign wire_6 = wire_6_0|wire_6_1;
  wire [7:0] wire_7;
  wire [7:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [7:0] wire_10_0;
  wire [7:0] wire_10_1;
  assign wire_10 = wire_10_0|wire_10_1;
  wire [0:0] wire_11;
  wire [7:0] wire_12;
  wire [7:0] wire_13;
  wire [7:0] wire_14;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  wire [0:0] wire_17;
  wire [7:0] wire_18;
  wire [7:0] wire_19;
  wire [0:0] wire_20;
  wire [7:0] wire_21;
  wire [7:0] wire_21_0;
  wire [7:0] wire_21_1;
  assign wire_21 = wire_21_0|wire_21_1;
  wire [7:0] wire_22;
  wire [7:0] wire_22_0;
  wire [7:0] wire_22_1;
  assign wire_22 = wire_22_0|wire_22_1;
  wire [0:0] wire_23;
  wire [7:0] wire_24;
  wire [7:0] wire_24_0;
  wire [7:0] wire_24_1;
  assign wire_24 = wire_24_0|wire_24_1;
  wire [7:0] wire_25;
  wire [0:0] wire_26;
  wire [7:0] wire_27;
  wire [7:0] wire_28;
  wire [7:0] wire_29;
  wire [7:0] wire_30;
  wire [7:0] wire_30_0;
  wire [7:0] wire_30_1;
  assign wire_30 = wire_30_0|wire_30_1;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [63:0] wire_33;
  assign wire_33 = Input;
  wire [7:0] wire_34;
  wire [7:0] wire_35;
  wire [7:0] wire_35_0;
  wire [7:0] wire_35_1;
  assign wire_35 = wire_35_0|wire_35_1;
  assign Output = wire_35;
  wire [7:0] wire_36;
  wire [7:0] wire_36_0;
  wire [7:0] wire_36_1;
  assign wire_36 = wire_36_0|wire_36_1;
  wire [7:0] wire_37;
  wire [7:0] wire_38;
  wire [7:0] wire_39;
  wire [0:0] wire_40;
  wire [7:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [7:0] wire_48;

endmodule
