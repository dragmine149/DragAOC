module Day2Part2z_Noz_Clean (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_Constant # (.UUID(64'd1726993617052590723 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFFFFFFFFFFFFFFFF)) Constant64_0 (.out(wire_56));
  TC_FileLoader # (.UUID(64'd3987767967543158583 ^ UUID), .DEFAULT_FILE_NAME("day2_modified")) FileLoader_1 (.clk(clk), .rst(rst), .en(wire_71), .address(wire_35), .out(wire_63_0));
  TC_Constant # (.UUID(64'd337803116546834142 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_2 (.out(wire_71));
  TC_LessU # (.UUID(64'd2415299641673726094 ^ UUID), .BIT_WIDTH(64'd64)) LessU64_3 (.in0(wire_90), .in1(wire_35), .out(wire_32));
  TC_FileLoader # (.UUID(64'd4235385288069024156 ^ UUID), .DEFAULT_FILE_NAME("day2_test_1")) FileLoader_4 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_35), .out(wire_63_1));
  TC_Constant # (.UUID(64'd1484234401691717814 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_5 (.out());
  TC_DelayLine # (.UUID(64'd2141883989358176841 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_6 (.clk(clk), .rst(rst), .in(wire_79), .out(wire_5));
  TC_Add # (.UUID(64'd3665390526026043059 ^ UUID), .BIT_WIDTH(64'd64)) Add64_7 (.in0({{56{1'b0}}, wire_28 }), .in1(wire_35), .ci(1'd0), .out(wire_61), .co());
  TC_Counter # (.UUID(64'd3781882184507484018 ^ UUID), .BIT_WIDTH(64'd64), .count(64'd1)) Counter64_8 (.clk(clk), .rst(rst), .save(wire_38), .in(wire_19), .out(wire_11));
  TC_Not # (.UUID(64'd2915069602117248147 ^ UUID), .BIT_WIDTH(64'd1)) Not_9 (.in(wire_32), .out(wire_66));
  TC_And # (.UUID(64'd4444366698480428793 ^ UUID), .BIT_WIDTH(64'd1)) And_10 (.in0(wire_9), .in1(wire_32), .out(wire_34));
  TC_Or # (.UUID(64'd1455535717111312185 ^ UUID), .BIT_WIDTH(64'd1)) Or_11 (.in0(wire_55), .in1(wire_34), .out(wire_38));
  TC_Not # (.UUID(64'd4292279915901693506 ^ UUID), .BIT_WIDTH(64'd1)) Not_12 (.in(wire_9), .out(wire_55));
  TC_Switch # (.UUID(64'd259253643073170517 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_13 (.en(wire_66), .in(wire_11), .out(wire_2_1));
  TC_Counter # (.UUID(64'd4027361701724138616 ^ UUID), .BIT_WIDTH(64'd64), .count(64'd1)) Counter64_14 (.clk(clk), .rst(rst), .save(wire_46), .in(wire_43), .out(wire_14));
  TC_Ram # (.UUID(64'd3231836939472590219 ^ UUID), .WORD_WIDTH(64'd64), .WORD_COUNT(64'd1250)) Ram_15 (.clk(clk), .rst(rst), .load(wire_12), .save(wire_20), .address(wire_2[31:0]), .in0(wire_1), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_23), .out1(), .out2(), .out3());
  TC_Halt # (.UUID(64'd1646709671390234641 ^ UUID), .HALT_MESSAGE("Program finished!")) Halt_16 (.clk(clk), .rst(rst), .en(wire_68));
  TC_NoteSound # (.UUID(64'd2856162216424263791 ^ UUID)) NoteSound_17 (.clk(clk), .rst(rst), .command({{7{1'b0}}, wire_68 }), .note(wire_86), .pitch(8'd0));
  TC_Constant # (.UUID(64'd3448097267265053438 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h28)) Constant8_18 (.out(wire_86));
  TC_Not # (.UUID(64'd1023328388184503186 ^ UUID), .BIT_WIDTH(64'd1)) Not_19 (.in(wire_34), .out(wire_53));
  TC_DelayLine # (.UUID(64'd4092965687359902133 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_20 (.clk(clk), .rst(rst), .in(wire_27), .out(wire_80));
  TC_Mux # (.UUID(64'd316725708318265243 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_21 (.sel(wire_9), .in0(wire_56), .in1(wire_80), .out(wire_35));
  TC_Switch # (.UUID(64'd3903258603175327041 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_22 (.en(wire_65), .in(wire_23), .out(wire_6));
  TC_Switch # (.UUID(64'd1710097796709442780 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_23 (.en(wire_18), .in(wire_23), .out(wire_15));
  TC_Switch # (.UUID(64'd3052143593441878759 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_24 (.en(wire_4), .in(wire_26), .out(wire_2_3));
  TC_Constant # (.UUID(64'd3240501465042579115 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_25 (.out(wire_85));
  TC_Not # (.UUID(64'd1867582932362601439 ^ UUID), .BIT_WIDTH(64'd1)) Not_26 (.in(wire_46), .out(wire_49));
  TC_DelayLine # (.UUID(64'd2677504830674658084 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_27 (.clk(clk), .rst(rst), .in(wire_0), .out(wire_51));
  TC_Switch # (.UUID(64'd1725179244806057793 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_28 (.en(wire_60), .in(wire_6), .out(wire_0));
  TC_DelayLine # (.UUID(64'd1784992797701007900 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_29 (.clk(clk), .rst(rst), .in(wire_60), .out(wire_25));
  TC_DelayLine # (.UUID(64'd4350311000933170162 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_30 (.clk(clk), .rst(rst), .in(wire_18), .out(wire_36));
  TC_Switch # (.UUID(64'd4182440545682965520 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_31 (.en(wire_70), .in(wire_15), .out(wire_47));
  TC_DelayLine # (.UUID(64'd247377800554737393 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_32 (.clk(clk), .rst(rst), .in(wire_47), .out(wire_81));
  TC_DelayLine # (.UUID(64'd3700638478856170501 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_33 (.clk(clk), .rst(rst), .in(wire_70), .out(wire_87));
  TC_Switch # (.UUID(64'd3804153078929315197 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_34 (.en(wire_25), .in(wire_51), .out(wire_26_0));
  TC_Switch # (.UUID(64'd79719301686403854 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_35 (.en(wire_87), .in(wire_81), .out(wire_26_1));
  TC_Add # (.UUID(64'd1069550484725226130 ^ UUID), .BIT_WIDTH(64'd64)) Add64_36 (.in0(wire_16), .in1(wire_59), .ci(1'd0), .out(wire_94), .co());
  TC_Mul # (.UUID(64'd924182476717345043 ^ UUID), .BIT_WIDTH(64'd64)) Mul64_37 (.in0(wire_16), .in1(wire_59), .out0(wire_96), .out1());
  TC_Switch # (.UUID(64'd935510424511562668 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_38 (.en(wire_39), .in(wire_94), .out(wire_7_1));
  TC_Switch # (.UUID(64'd3389748284807452395 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_39 (.en(wire_58), .in(wire_96), .out(wire_7_0));
  TC_Halt # (.UUID(64'd3795677300099293191 ^ UUID), .HALT_MESSAGE("Opcode 99 Reached!")) Halt_40 (.clk(clk), .rst(rst), .en(1'd0));
  TC_Switch # (.UUID(64'd1224855048361981157 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_41 (.en(wire_33), .in(wire_7), .out(wire_1_0));
  TC_And # (.UUID(64'd4423175184107256786 ^ UUID), .BIT_WIDTH(64'd1)) And_42 (.in0(wire_50), .in1(wire_82), .out(wire_33));
  TC_Constant # (.UUID(64'd2201783711648500038 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_43 (.out(wire_82));
  TC_Not # (.UUID(64'd3940936562307563579 ^ UUID), .BIT_WIDTH(64'd1)) Not_44 (.in(wire_33), .out(wire_74));
  TC_DelayLine # (.UUID(64'd366563469061908473 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_45 (.clk(clk), .rst(rst), .in(wire_74), .out(wire_44));
  TC_Not # (.UUID(64'd23546066323564917 ^ UUID), .BIT_WIDTH(64'd1)) Not_46 (.in(wire_34), .out(wire_41));
  TC_Or3 # (.UUID(64'd1565632499214780517 ^ UUID), .BIT_WIDTH(64'd1)) Or3_47 (.in0(wire_3), .in1(wire_21), .in2(wire_53), .out(wire_46_1));
  TC_Not # (.UUID(64'd601742535760828746 ^ UUID), .BIT_WIDTH(64'd1)) Not_48 (.in(wire_54), .out(wire_24));
  TC_DelayLine # (.UUID(64'd1263282884327671549 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_49 (.clk(clk), .rst(rst), .in(wire_65), .out(wire_13));
  TC_Not # (.UUID(64'd4567426784455268513 ^ UUID), .BIT_WIDTH(64'd1)) Not_50 (.in(wire_13), .out(wire_77));
  TC_Not # (.UUID(64'd4522425577002129070 ^ UUID), .BIT_WIDTH(64'd1)) Not_51 (.in(wire_36), .out(wire_69));
  TC_Or # (.UUID(64'd571059853550174113 ^ UUID), .BIT_WIDTH(64'd1)) Or_52 (.in0(wire_37), .in1(wire_33), .out(wire_21));
  TC_FileLoader # (.UUID(64'd4032583951989155851 ^ UUID), .DEFAULT_FILE_NAME("day2_test_2")) FileLoader_53 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_35), .out(wire_63_2));
  TC_Constant # (.UUID(64'd1883781277529937826 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_54 (.out());
  TC_Constant # (.UUID(64'd4566527038733230091 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_55 (.out());
  TC_Constant # (.UUID(64'd3138890809031518109 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_56 (.out());
  TC_Constant # (.UUID(64'd2829021048917779791 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_57 (.out());
  TC_Constant # (.UUID(64'd1405985673201260239 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_58 (.out());
  TC_Constant # (.UUID(64'd3716163551666950261 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_59 (.out());
  TC_Constant # (.UUID(64'd4023943151529497828 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_60 (.out());
  TC_Constant # (.UUID(64'd2532988701438288488 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_61 (.out());
  TC_Constant # (.UUID(64'd4214058095318520776 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_62 (.out());
  TC_Constant # (.UUID(64'd958940107339709111 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_63 (.out());
  TC_Constant # (.UUID(64'd2113422115012713154 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_64 (.out());
  TC_Constant # (.UUID(64'd372203303927728035 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_65 (.out());
  TC_Constant # (.UUID(64'd4215445727210423365 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_66 (.out());
  TC_Constant # (.UUID(64'd4177145269316879433 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_67 (.out());
  TC_FileLoader # (.UUID(64'd3305349617174586722 ^ UUID), .DEFAULT_FILE_NAME("day2_test_3")) FileLoader_68 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_35), .out(wire_63_3));
  TC_FileLoader # (.UUID(64'd231382507668522051 ^ UUID), .DEFAULT_FILE_NAME("day2_test_4")) FileLoader_69 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_35), .out(wire_63_4));
  TC_FileLoader # (.UUID(64'd1231532553883646540 ^ UUID), .DEFAULT_FILE_NAME("day2_test_5")) FileLoader_70 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_35), .out(wire_63_5));
  TC_Equal # (.UUID(64'd2821604189245118802 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_71 (.in0(wire_11), .in1({{56{1'b0}}, wire_84 }), .out(wire_10));
  TC_Equal # (.UUID(64'd834176164977634459 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_72 (.in0(wire_11), .in1({{56{1'b0}}, wire_62 }), .out(wire_8));
  TC_Constant # (.UUID(64'd1065572658605867570 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_73 (.out(wire_84));
  TC_Constant # (.UUID(64'd991865579609327770 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_74 (.out(wire_62));
  TC_Switch # (.UUID(64'd1746571703522486786 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_75 (.en(wire_10), .in(wire_95), .out(wire_57_0));
  TC_Switch # (.UUID(64'd1454525939490593477 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_76 (.en(wire_8), .in(wire_93), .out(wire_57_1));
  TC_Switch # (.UUID(64'd1728873000476622687 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_77 (.en(wire_29), .in(wire_72[7:0]), .out(wire_57_2));
  TC_Nor # (.UUID(64'd4535549015773012659 ^ UUID), .BIT_WIDTH(64'd1)) Nor_78 (.in0(wire_10), .in1(wire_8), .out(wire_29));
  TC_Equal # (.UUID(64'd4382296156982196310 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_79 (.in0(wire_23), .in1(wire_64), .out(wire_45));
  TC_And # (.UUID(64'd1888702582889417503 ^ UUID), .BIT_WIDTH(64'd1)) And_80 (.in0(wire_45), .in1(wire_37), .out(wire_17));
  TC_Halt # (.UUID(64'd4563628704689697466 ^ UUID), .HALT_MESSAGE("Number pair found!")) Halt_81 (.clk(clk), .rst(rst), .en(wire_17));
  TC_Constant # (.UUID(64'd2825119468061589370 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h12C74E0)) Constant64_82 (.out(wire_64));
  TC_Switch # (.UUID(64'd2786939255044915453 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_83 (.en(wire_31), .in(wire_11), .out(wire_19));
  TC_Halt # (.UUID(64'd173880931492206516 ^ UUID), .HALT_MESSAGE("Memory Cleared")) Halt_84 (.clk(clk), .rst(rst), .en(1'd0));
  TC_And # (.UUID(64'd1254581417745991036 ^ UUID), .BIT_WIDTH(64'd1)) And_85 (.in0(wire_37), .in1(wire_75), .out(wire_22));
  TC_Switch # (.UUID(64'd2236419431862390674 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_86 (.en(wire_31), .in(wire_61), .out(wire_27));
  TC_Not # (.UUID(64'd895591967131792673 ^ UUID), .BIT_WIDTH(64'd1)) Not_87 (.in(wire_22), .out(wire_31));
  TC_Switch # (.UUID(64'd1341671548569791167 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_88 (.en(wire_67), .in(wire_14), .out(wire_43));
  TC_Not # (.UUID(64'd1026398734405901705 ^ UUID), .BIT_WIDTH(64'd1)) Not_89 (.in(wire_67), .out(wire_91));
  TC_DelayLine # (.UUID(64'd3662433804087744831 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_90 (.clk(clk), .rst(rst), .in(wire_31), .out(wire_67));
  TC_Halt # (.UUID(64'd2336335384836364761 ^ UUID), .HALT_MESSAGE("Panic! Not found number within time frame!")) Halt_91 (.clk(clk), .rst(rst), .en(wire_76));
  QuickSave # (.UUID(64'd2695330121804011308 ^ UUID)) QuickSave_92 (.clk(clk), .rst(rst), .Value(wire_63), .\Number_(stored) (wire_90), .\Saved?_1 (wire_9), .\Saved?_2 ());
  BytesToNumbersz_3 # (.UUID(64'd1729469431074511873 ^ UUID)) BytesToNumbersz_3_93 (.clk(clk), .rst(rst), .Main_8b(wire_63), .Carry_In(wire_5), .Output(wire_79), .Offset(wire_28), .Value(wire_72));
  OnOrOff # (.UUID(64'd3163142382288365090 ^ UUID)) OnOrOff_94 (.clk(clk), .rst(rst), .Input(wire_66), .Output(wire_20_1));
  flippedzm64bzmswitch # (.UUID(64'd2031059029553199162 ^ UUID)) flippedzm64bzmswitch_95 (.clk(clk), .rst(rst), .Input_1(wire_14), .Input_2(wire_49), .Output(wire_2_2));
  OnOrOff # (.UUID(64'd150349705086353648 ^ UUID)) OnOrOff_96 (.clk(clk), .rst(rst), .Input(wire_49), .Output(wire_12_1));
  OnOrOff # (.UUID(64'd224193335304047014 ^ UUID)) OnOrOff_97 (.clk(clk), .rst(rst), .Input(wire_83), .Output(wire_12_0));
  mand # (.UUID(64'd3349436745291189726 ^ UUID)) mand_98 (.clk(clk), .rst(rst), .Input_1(wire_3), .Input_2(wire_85), .Output(wire_83));
  mand # (.UUID(64'd242248694494001734 ^ UUID)) mand_99 (.clk(clk), .rst(rst), .Input_1(wire_34), .Input_2(wire_44), .Output(wire_54));
  flippedzm64bzmswitch # (.UUID(64'd1881707450118815654 ^ UUID)) flippedzm64bzmswitch_100 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_13), .Output(wire_78));
  OnOrOff # (.UUID(64'd4158355321388927517 ^ UUID)) OnOrOff_101 (.clk(clk), .rst(rst), .Input(wire_25), .Output(wire_3_0));
  flippedzm64bzmswitch # (.UUID(64'd558922318308219109 ^ UUID)) flippedzm64bzmswitch_102 (.clk(clk), .rst(rst), .Input_1(wire_15), .Input_2(wire_36), .Output(wire_88));
  OnOrOff # (.UUID(64'd3868852299644989347 ^ UUID)) OnOrOff_103 (.clk(clk), .rst(rst), .Input(wire_87), .Output(wire_3_1));
  Opcodez_zmz_1z_2z_99 # (.UUID(64'd1253066027045582023 ^ UUID)) Opcodez_zmz_1z_2z_99_104 (.clk(clk), .rst(rst), .Opcode(wire_42[7:0]), .Add(wire_39), .divide(wire_58), .halt(wire_37));
  OnOrOff # (.UUID(64'd779081389060044986 ^ UUID)) OnOrOff_105 (.clk(clk), .rst(rst), .Input(wire_33), .Output(wire_20_0));
  flippedzm64bzmswitch # (.UUID(64'd3330710435434371616 ^ UUID)) flippedzm64bzmswitch_106 (.clk(clk), .rst(rst), .Input_1(wire_40), .Input_2(wire_33), .Output(wire_2_0));
  flippedzm64bzmswitch # (.UUID(64'd3395453474976780481 ^ UUID)) flippedzm64bzmswitch_107 (.clk(clk), .rst(rst), .Input_1({{56{1'b0}}, wire_57 }), .Input_2(wire_41), .Output(wire_1_1));
  CellWritter # (.UUID(64'd1760994904368207804 ^ UUID)) CellWritter_108 (.clk(clk), .rst(rst), .Clear(wire_24), .Write(wire_12), .Value_1(wire_23), .Value_2(wire_42), .Written(wire_92));
  CellWritter # (.UUID(64'd2225673571882546958 ^ UUID)) CellWritter_109 (.clk(clk), .rst(rst), .Clear(wire_24), .Write(wire_13), .Value_1(wire_78), .Value_2(wire_16), .Written(wire_73));
  CellWritter # (.UUID(64'd640733034693975124 ^ UUID)) CellWritter_110 (.clk(clk), .rst(rst), .Clear(wire_24), .Write(wire_36), .Value_1(wire_88), .Value_2(wire_59), .Written(wire_52));
  mand # (.UUID(64'd2253745888330672149 ^ UUID)) mand_111 (.clk(clk), .rst(rst), .Input_1(wire_65), .Input_2(wire_77), .Output(wire_60));
  mand # (.UUID(64'd4089700112481536660 ^ UUID)) mand_112 (.clk(clk), .rst(rst), .Input_1(wire_18), .Input_2(wire_69), .Output(wire_70));
  CellWritter # (.UUID(64'd3735606448599014512 ^ UUID)) CellWritter_113 (.clk(clk), .rst(rst), .Clear(wire_24), .Write(wire_30), .Value_1(wire_23), .Value_2(wire_40), .Written(wire_50));
  mand # (.UUID(64'd1207172339067544539 ^ UUID)) mand_114 (.clk(clk), .rst(rst), .Input_1(wire_92), .Input_2(wire_12), .Output(wire_65));
  mand # (.UUID(64'd1055636189021926738 ^ UUID)) mand_115 (.clk(clk), .rst(rst), .Input_1(wire_73), .Input_2(wire_12), .Output(wire_18));
  mand # (.UUID(64'd3603338431621519469 ^ UUID)) mand_116 (.clk(clk), .rst(rst), .Input_1(wire_52), .Input_2(wire_12), .Output(wire_30));
  OnOrOff # (.UUID(64'd2326604957341175433 ^ UUID)) OnOrOff_117 (.clk(clk), .rst(rst), .Input(wire_37), .Output(wire_12_2));
  _99z_Counterz_Manual # (.UUID(64'd1622372112810930977 ^ UUID)) _99z_Counterz_Manual_118 (.clk(clk), .rst(rst), .Manual_Incrment(wire_89), .Out(wire_93), .Increment(wire_76));
  _99z_Counterz_Manual # (.UUID(64'd436698719286378264 ^ UUID)) _99z_Counterz_Manual_119 (.clk(clk), .rst(rst), .Manual_Incrment(wire_22), .Out(wire_95), .Increment(wire_89));
  _64zmany # (.UUID(64'd1931968964033189129 ^ UUID)) _64zmany_120 (.clk(clk), .rst(rst), .Input(wire_11), .Output(wire_75));
  OnOrOff # (.UUID(64'd4135007685282140821 ^ UUID)) OnOrOff_121 (.clk(clk), .rst(rst), .Input(wire_91), .Output(wire_46_0));
  TC_And # (.UUID(64'd166281153331008272 ^ UUID), .BIT_WIDTH(64'd1)) And_122 (.in0(wire_3), .in1(wire_48), .out(wire_4));
  TC_Not # (.UUID(64'd141376591780260008 ^ UUID), .BIT_WIDTH(64'd1)) Not_123 (.in(wire_37), .out(wire_48));

  wire [63:0] wire_0;
  wire [63:0] wire_1;
  wire [63:0] wire_1_0;
  wire [63:0] wire_1_1;
  assign wire_1 = wire_1_0|wire_1_1;
  wire [63:0] wire_2;
  wire [63:0] wire_2_0;
  wire [63:0] wire_2_1;
  wire [63:0] wire_2_2;
  wire [63:0] wire_2_3;
  assign wire_2 = wire_2_0|wire_2_1|wire_2_2|wire_2_3;
  wire [0:0] wire_3;
  wire [0:0] wire_3_0;
  wire [0:0] wire_3_1;
  assign wire_3 = wire_3_0|wire_3_1;
  wire [0:0] wire_4;
  wire [63:0] wire_5;
  wire [63:0] wire_6;
  wire [63:0] wire_7;
  wire [63:0] wire_7_0;
  wire [63:0] wire_7_1;
  assign wire_7 = wire_7_0|wire_7_1;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [63:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_12_0;
  wire [0:0] wire_12_1;
  wire [0:0] wire_12_2;
  assign wire_12 = wire_12_0|wire_12_1|wire_12_2;
  wire [0:0] wire_13;
  wire [63:0] wire_14;
  wire [63:0] wire_15;
  wire [63:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [63:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_20_0;
  wire [0:0] wire_20_1;
  assign wire_20 = wire_20_0|wire_20_1;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [63:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [63:0] wire_26;
  wire [63:0] wire_26_0;
  wire [63:0] wire_26_1;
  assign wire_26 = wire_26_0|wire_26_1;
  wire [63:0] wire_27;
  wire [7:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [63:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [63:0] wire_40;
  wire [0:0] wire_41;
  wire [63:0] wire_42;
  wire [63:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_46_0;
  wire [0:0] wire_46_1;
  assign wire_46 = wire_46_0|wire_46_1;
  wire [63:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [63:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [63:0] wire_56;
  wire [7:0] wire_57;
  wire [7:0] wire_57_0;
  wire [7:0] wire_57_1;
  wire [7:0] wire_57_2;
  assign wire_57 = wire_57_0|wire_57_1|wire_57_2;
  wire [0:0] wire_58;
  wire [63:0] wire_59;
  wire [0:0] wire_60;
  wire [63:0] wire_61;
  wire [7:0] wire_62;
  wire [63:0] wire_63;
  wire [63:0] wire_63_0;
  wire [63:0] wire_63_1;
  wire [63:0] wire_63_2;
  wire [63:0] wire_63_3;
  wire [63:0] wire_63_4;
  wire [63:0] wire_63_5;
  assign wire_63 = wire_63_0|wire_63_1|wire_63_2|wire_63_3|wire_63_4|wire_63_5;
  wire [63:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  assign wire_68 = 0;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [63:0] wire_72;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [63:0] wire_78;
  wire [63:0] wire_79;
  wire [63:0] wire_80;
  wire [63:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [7:0] wire_84;
  wire [0:0] wire_85;
  wire [7:0] wire_86;
  wire [0:0] wire_87;
  wire [63:0] wire_88;
  wire [0:0] wire_89;
  wire [63:0] wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  wire [7:0] wire_93;
  wire [63:0] wire_94;
  wire [7:0] wire_95;
  wire [63:0] wire_96;

endmodule
