module is0z_32b (clk, rst, Input, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [31:0] Input;
  output  wire [0:0] Output;

  TC_Splitter32 # (.UUID(64'd3807558696634726507 ^ UUID)) Splitter32_0 (.in(wire_4), .out0(wire_9), .out1(wire_5), .out2(wire_1), .out3(wire_2));
  TC_Maker16 # (.UUID(64'd4058533878944925470 ^ UUID)) Maker16_1 (.in0(wire_9), .in1(wire_5), .out(wire_7));
  TC_Maker16 # (.UUID(64'd1600105428663763521 ^ UUID)) Maker16_2 (.in0(wire_1), .in1(wire_2), .out(wire_3));
  is0 # (.UUID(64'd56137896704869034 ^ UUID)) is0_3 (.clk(clk), .rst(rst), .Input(wire_7), .Output(wire_0));
  is0 # (.UUID(64'd1173233436144774023 ^ UUID)) is0_4 (.clk(clk), .rst(rst), .Input(wire_3), .Output(wire_8));
  TC_And # (.UUID(64'd3554763759628229062 ^ UUID), .BIT_WIDTH(64'd1)) And_5 (.in0(wire_0), .in1(wire_8), .out(wire_6));

  wire [0:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_2;
  wire [15:0] wire_3;
  wire [31:0] wire_4;
  assign wire_4 = Input;
  wire [7:0] wire_5;
  wire [0:0] wire_6;
  assign Output = wire_6;
  wire [15:0] wire_7;
  wire [0:0] wire_8;
  wire [7:0] wire_9;

endmodule
