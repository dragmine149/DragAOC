module Day4Part1z_2 (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_FileLoader # (.UUID(64'd1300333077211007914 ^ UUID), .DEFAULT_FILE_NAME("day4")) FileLoader_0 (.clk(clk), .rst(rst), .en(wire_60), .address({{56{1'b0}}, wire_39 }), .out(wire_16));
  TC_Constant # (.UUID(64'd614705877810942359 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_1 (.out(wire_60));
  TC_IndexerByte # (.UUID(64'd3259875342327518678 ^ UUID), .INDEX(64'd0)) IndexerByte_2 (.in(wire_16), .out(wire_25));
  TC_Constant # (.UUID(64'd2881157116684703501 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_3 (.out(wire_33));
  TC_IndexerByte # (.UUID(64'd3282167999629572026 ^ UUID), .INDEX(64'd0)) IndexerByte_4 (.in(wire_4), .out(wire_10));
  TC_IndexerByte # (.UUID(64'd344938491191684993 ^ UUID), .INDEX(64'd1)) IndexerByte_5 (.in(wire_4), .out(wire_52));
  TC_IndexerByte # (.UUID(64'd3057145202194435591 ^ UUID), .INDEX(64'd2)) IndexerByte_6 (.in(wire_4), .out(wire_54));
  TC_IndexerByte # (.UUID(64'd196694779505405906 ^ UUID), .INDEX(64'd3)) IndexerByte_7 (.in(wire_4), .out(wire_37));
  TC_IndexerByte # (.UUID(64'd195480252778983173 ^ UUID), .INDEX(64'd4)) IndexerByte_8 (.in(wire_4), .out(wire_31));
  TC_IndexerByte # (.UUID(64'd2249681588834216334 ^ UUID), .INDEX(64'd5)) IndexerByte_9 (.in(wire_4), .out(wire_9));
  TC_Maker64 # (.UUID(64'd2041678736802242094 ^ UUID)) Maker64_10 (.in0(wire_58), .in1(wire_56), .in2(wire_27), .in3(wire_44), .in4(wire_2), .in5(wire_74), .in6(8'd0), .in7(8'd0), .out(wire_4));
  TC_DelayLine # (.UUID(64'd1478884666127726678 ^ UUID), .BIT_WIDTH(64'd8)) DelayLine8_11 (.clk(clk), .rst(rst), .in(wire_34), .out(wire_39));
  TC_Constant # (.UUID(64'd4230246302748610089 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_12 (.out(wire_34));
  TC_IndexerByte # (.UUID(64'd3885874403913997322 ^ UUID), .INDEX(64'd1)) IndexerByte_13 (.in(wire_16), .out(wire_71));
  TC_IndexerByte # (.UUID(64'd2749811280805536878 ^ UUID), .INDEX(64'd2)) IndexerByte_14 (.in(wire_16), .out(wire_38));
  TC_IndexerByte # (.UUID(64'd3113000412030619556 ^ UUID), .INDEX(64'd3)) IndexerByte_15 (.in(wire_16), .out(wire_59));
  TC_IndexerByte # (.UUID(64'd3058128748266773168 ^ UUID), .INDEX(64'd4)) IndexerByte_16 (.in(wire_16), .out(wire_13));
  TC_IndexerByte # (.UUID(64'd3726479596336349432 ^ UUID), .INDEX(64'd5)) IndexerByte_17 (.in(wire_16), .out(wire_67));
  TC_Splitter64 # (.UUID(64'd1715894660434795144 ^ UUID)) Splitter64_18 (.in(wire_51), .out0(wire_43), .out1(wire_0), .out2(wire_53), .out3(wire_26), .out4(wire_48), .out5(wire_21), .out6(), .out7());
  TC_Switch # (.UUID(64'd3083524623901623221 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_19 (.en(wire_23), .in(wire_4), .out(wire_51));
  TC_Not # (.UUID(64'd1741588675539327596 ^ UUID), .BIT_WIDTH(64'd1)) Not_20 (.in(wire_15), .out(wire_23));
  TC_Counter # (.UUID(64'd2796646339049657840 ^ UUID), .BIT_WIDTH(64'd16), .count(16'd1)) Counter16_21 (.clk(clk), .rst(rst), .save(wire_57), .in(wire_8), .out(wire_8));
  TC_Not # (.UUID(64'd262671911581901502 ^ UUID), .BIT_WIDTH(64'd1)) Not_22 (.in(wire_73), .out(wire_57));
  TC_Halt # (.UUID(64'd2373505150995397943 ^ UUID), .HALT_MESSAGE("Upper limit reached")) Halt_23 (.clk(clk), .rst(rst), .en(wire_70));
  TC_Switch # (.UUID(64'd4386075278005230458 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_24 (.en(wire_23), .in(wire_45), .out(wire_70));
  TC_LessI # (.UUID(64'd3292654551045928704 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_25 (.in0(wire_3), .in1(wire_1), .out(wire_29));
  TC_LessI # (.UUID(64'd3747362352843898306 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_26 (.in0(wire_5), .in1(wire_3), .out(wire_55));
  TC_LessI # (.UUID(64'd4227878923150009143 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_27 (.in0(wire_14), .in1(wire_5), .out(wire_65));
  TC_LessI # (.UUID(64'd4090912352078921077 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_28 (.in0(wire_28), .in1(wire_14), .out(wire_63));
  TC_LessI # (.UUID(64'd2040532423834977934 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_29 (.in0(wire_50), .in1(wire_28), .out(wire_69));
  TC_Not # (.UUID(64'd366707461536672635 ^ UUID), .BIT_WIDTH(64'd1)) Not_30 (.in(wire_69), .out(wire_30));
  TC_Not # (.UUID(64'd2939040142042526066 ^ UUID), .BIT_WIDTH(64'd1)) Not_31 (.in(wire_63), .out(wire_41));
  TC_Not # (.UUID(64'd1398917821098271411 ^ UUID), .BIT_WIDTH(64'd1)) Not_32 (.in(wire_65), .out(wire_72));
  TC_Not # (.UUID(64'd3712273125459795596 ^ UUID), .BIT_WIDTH(64'd1)) Not_33 (.in(wire_55), .out(wire_47));
  TC_Not # (.UUID(64'd349618724439403530 ^ UUID), .BIT_WIDTH(64'd1)) Not_34 (.in(wire_29), .out(wire_40));
  TC_And # (.UUID(64'd949179814438959664 ^ UUID), .BIT_WIDTH(64'd1)) And_35 (.in0(wire_20), .in1(wire_18), .out(wire_64));
  TC_Switch # (.UUID(64'd3806424035603758608 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_36 (.en(wire_23), .in(wire_64), .out(wire_73));
  NotTick # (.UUID(64'd988254291887862844 ^ UUID)) NotTick_37 (.clk(clk), .rst(rst), .Output(wire_15));
  ByteToNumber # (.UUID(64'd2290549341218488923 ^ UUID)) ByteToNumber_38 (.clk(clk), .rst(rst), .Input(wire_25), .Output(wire_58));
  ByteToNumber # (.UUID(64'd4267877789773175085 ^ UUID)) ByteToNumber_39 (.clk(clk), .rst(rst), .Input(wire_71), .Output(wire_56));
  ByteToNumber # (.UUID(64'd803095588841364073 ^ UUID)) ByteToNumber_40 (.clk(clk), .rst(rst), .Input(wire_38), .Output(wire_27));
  ByteToNumber # (.UUID(64'd677672594194363867 ^ UUID)) ByteToNumber_41 (.clk(clk), .rst(rst), .Input(wire_59), .Output(wire_44));
  ByteToNumber # (.UUID(64'd2617233141476735101 ^ UUID)) ByteToNumber_42 (.clk(clk), .rst(rst), .Input(wire_13), .Output(wire_2));
  ByteToNumber # (.UUID(64'd3235338507986847377 ^ UUID)) ByteToNumber_43 (.clk(clk), .rst(rst), .Input(wire_67), .Output(wire_74));
  _4beq # (.UUID(64'd4084947534873581742 ^ UUID)) _4beq_44 (.clk(clk), .rst(rst), .Input_1(wire_1), .Input_2(wire_3), .Output(wire_36));
  _4beq # (.UUID(64'd837930388802506938 ^ UUID)) _4beq_45 (.clk(clk), .rst(rst), .Input_1(wire_3), .Input_2(wire_5), .Output(wire_62));
  _4beq # (.UUID(64'd1001160964423906324 ^ UUID)) _4beq_46 (.clk(clk), .rst(rst), .Input_1(wire_5), .Input_2(wire_14), .Output(wire_7));
  _4beq # (.UUID(64'd4024915304172217312 ^ UUID)) _4beq_47 (.clk(clk), .rst(rst), .Input_1(wire_14), .Input_2(wire_28), .Output(wire_11));
  _4beq # (.UUID(64'd3801586074555563384 ^ UUID)) _4beq_48 (.clk(clk), .rst(rst), .Input_1(wire_28), .Input_2(wire_50), .Output(wire_75));
  OnOrOff # (.UUID(64'd2794213930716429597 ^ UUID)) OnOrOff_49 (.clk(clk), .rst(rst), .Input(wire_62), .Output(wire_20_0));
  OnOrOff # (.UUID(64'd321309780266364927 ^ UUID)) OnOrOff_50 (.clk(clk), .rst(rst), .Input(wire_7), .Output(wire_20_2));
  OnOrOff # (.UUID(64'd2791637861636592922 ^ UUID)) OnOrOff_51 (.clk(clk), .rst(rst), .Input(wire_11), .Output(wire_20_3));
  OnOrOff # (.UUID(64'd4363176194552780331 ^ UUID)) OnOrOff_52 (.clk(clk), .rst(rst), .Input(wire_75), .Output(wire_20_4));
  OnOrOff # (.UUID(64'd2565202741671842960 ^ UUID)) OnOrOff_53 (.clk(clk), .rst(rst), .Input(wire_36), .Output(wire_20_1));
  mand # (.UUID(64'd2743742951316189243 ^ UUID)) mand_54 (.clk(clk), .rst(rst), .Input_1(wire_40), .Input_2(wire_47), .Output(wire_68));
  mand # (.UUID(64'd2942067753606735184 ^ UUID)) mand_55 (.clk(clk), .rst(rst), .Input_1(wire_72), .Input_2(wire_41), .Output(wire_6));
  mand # (.UUID(64'd18958839450887314 ^ UUID)) mand_56 (.clk(clk), .rst(rst), .Input_1(wire_68), .Input_2(wire_61), .Output(wire_18));
  mand # (.UUID(64'd3212422335951933954 ^ UUID)) mand_57 (.clk(clk), .rst(rst), .Input_1(wire_6), .Input_2(wire_30), .Output(wire_61));
  RangeChecker # (.UUID(64'd2690237951565181585 ^ UUID)) RangeChecker_58 (.clk(clk), .rst(rst), .Input_1(wire_0), .Input_2(wire_3), .Input_3(wire_43), .Input_4(wire_1), .Input_5(wire_21), .Input_6(wire_50), .Input_7(wire_48), .Input_8(wire_28), .Input_9(wire_26), .Input_10(wire_14), .Input_11(wire_53), .Input_12(wire_5), .Output(wire_45));
  Cellz_2 # (.UUID(64'd2681121728217391920 ^ UUID)) Cellz_2_59 (.clk(clk), .rst(rst), .Increment(wire_19), .Overwrite(wire_10), .Global_Overwrite(wire_15), .Previous(8'd0), .Output(wire_1), .Increment_Next());
  Cellz_2 # (.UUID(64'd3469695128675857344 ^ UUID)) Cellz_2_60 (.clk(clk), .rst(rst), .Increment(wire_35), .Overwrite(wire_52), .Global_Overwrite(wire_15), .Previous(wire_1), .Output(wire_3), .Increment_Next(wire_19));
  Cellz_2 # (.UUID(64'd2464365340593423882 ^ UUID)) Cellz_2_61 (.clk(clk), .rst(rst), .Increment(wire_32), .Overwrite(wire_54), .Global_Overwrite(wire_15), .Previous(wire_3), .Output(wire_5), .Increment_Next(wire_35));
  Cellz_2 # (.UUID(64'd403371948968645324 ^ UUID)) Cellz_2_62 (.clk(clk), .rst(rst), .Increment(wire_49), .Overwrite(wire_37), .Global_Overwrite(wire_15), .Previous(wire_5), .Output(wire_14), .Increment_Next(wire_32));
  Cellz_2 # (.UUID(64'd1534890721647203275 ^ UUID)) Cellz_2_63 (.clk(clk), .rst(rst), .Increment(wire_42), .Overwrite(wire_31), .Global_Overwrite(wire_15), .Previous(wire_14), .Output(wire_28), .Increment_Next(wire_49));
  Cellz_2 # (.UUID(64'd2165210612851354234 ^ UUID)) Cellz_2_64 (.clk(clk), .rst(rst), .Increment(wire_22), .Overwrite(wire_9), .Global_Overwrite(wire_15), .Previous(wire_28), .Output(wire_50), .Increment_Next(wire_42));
  TC_Switch # (.UUID(64'd3815757842053566393 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_65 (.en(wire_12), .in(wire_33), .out(wire_22));
  OnOrOff # (.UUID(64'd129879025491825736 ^ UUID)) OnOrOff_66 (.clk(clk), .rst(rst), .Input(wire_19), .Output(wire_24_0));
  OnOrOff # (.UUID(64'd2069905977387596 ^ UUID)) OnOrOff_67 (.clk(clk), .rst(rst), .Input(wire_35), .Output(wire_24_1));
  OnOrOff # (.UUID(64'd4020034695276023527 ^ UUID)) OnOrOff_68 (.clk(clk), .rst(rst), .Input(wire_32), .Output(wire_17_2));
  OnOrOff # (.UUID(64'd3681849683264036923 ^ UUID)) OnOrOff_69 (.clk(clk), .rst(rst), .Input(wire_49), .Output(wire_17_1));
  OnOrOff # (.UUID(64'd1477728482954482203 ^ UUID)) OnOrOff_70 (.clk(clk), .rst(rst), .Input(wire_42), .Output(wire_17_0));
  TC_Not # (.UUID(64'd4517909894909000332 ^ UUID), .BIT_WIDTH(64'd1)) Not_71 (.in(wire_66), .out(wire_12));
  TC_DelayLine # (.UUID(64'd1998668017909422993 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_72 (.clk(clk), .rst(rst), .in(wire_17), .out(wire_66));
  TC_DelayLine # (.UUID(64'd2142609526691430932 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_73 (.clk(clk), .rst(rst), .in(wire_24), .out(wire_46));
  OnOrOff # (.UUID(64'd2385286065099818749 ^ UUID)) OnOrOff_74 (.clk(clk), .rst(rst), .Input(wire_46), .Output(wire_17_3));

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_3;
  wire [63:0] wire_4;
  wire [7:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [15:0] wire_8;
  wire [7:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [7:0] wire_13;
  wire [7:0] wire_14;
  wire [0:0] wire_15;
  wire [63:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_17_0;
  wire [0:0] wire_17_1;
  wire [0:0] wire_17_2;
  wire [0:0] wire_17_3;
  assign wire_17 = wire_17_0|wire_17_1|wire_17_2|wire_17_3;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_20_0;
  wire [0:0] wire_20_1;
  wire [0:0] wire_20_2;
  wire [0:0] wire_20_3;
  wire [0:0] wire_20_4;
  assign wire_20 = wire_20_0|wire_20_1|wire_20_2|wire_20_3|wire_20_4;
  wire [7:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_24_0;
  wire [0:0] wire_24_1;
  assign wire_24 = wire_24_0|wire_24_1;
  wire [7:0] wire_25;
  wire [7:0] wire_26;
  wire [7:0] wire_27;
  wire [7:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [7:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [7:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [7:0] wire_37;
  wire [7:0] wire_38;
  wire [7:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [7:0] wire_43;
  wire [7:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [7:0] wire_48;
  wire [0:0] wire_49;
  wire [7:0] wire_50;
  wire [63:0] wire_51;
  wire [7:0] wire_52;
  wire [7:0] wire_53;
  wire [7:0] wire_54;
  wire [0:0] wire_55;
  wire [7:0] wire_56;
  wire [0:0] wire_57;
  wire [7:0] wire_58;
  wire [7:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [7:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [7:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [7:0] wire_74;
  wire [0:0] wire_75;

endmodule
