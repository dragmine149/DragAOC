module BytesToNumbersz_3 (clk, rst, Main_8b, Carry_In, Output, Offset, Value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [63:0] Main_8b;
  input  wire [63:0] Carry_In;
  output  wire [63:0] Output;
  output  wire [7:0] Offset;
  output  wire [63:0] Value;

  TC_Not # (.UUID(64'd409634758639379263 ^ UUID), .BIT_WIDTH(64'd1)) Not_0 (.in(wire_11), .out(wire_32));
  TC_Not # (.UUID(64'd1881815919858912192 ^ UUID), .BIT_WIDTH(64'd1)) Not_1 (.in(wire_53), .out(wire_28));
  TC_Not # (.UUID(64'd937236105432722860 ^ UUID), .BIT_WIDTH(64'd1)) Not_2 (.in(wire_6), .out(wire_5));
  TC_Not # (.UUID(64'd2594318732283820489 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_0), .out(wire_13));
  TC_Not # (.UUID(64'd174051712027247617 ^ UUID), .BIT_WIDTH(64'd1)) Not_4 (.in(wire_2), .out(wire_24));
  TC_Not # (.UUID(64'd181353414880786372 ^ UUID), .BIT_WIDTH(64'd1)) Not_5 (.in(wire_7), .out(wire_43));
  TC_Not # (.UUID(64'd4265371004147168272 ^ UUID), .BIT_WIDTH(64'd1)) Not_6 (.in(wire_12), .out(wire_50));
  TC_Not # (.UUID(64'd3630341913520932399 ^ UUID), .BIT_WIDTH(64'd1)) Not_7 (.in(wire_14), .out(wire_16));
  TC_Switch # (.UUID(64'd207939087145431957 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_8 (.en(wire_14), .in(wire_20), .out(wire_46));
  TC_Switch # (.UUID(64'd2304949746688299596 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_9 (.en(wire_12), .in(wire_54), .out(wire_71));
  TC_Switch # (.UUID(64'd1652140659488077705 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_10 (.en(wire_7), .in(wire_49), .out(wire_76));
  TC_Switch # (.UUID(64'd476386494605725266 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_11 (.en(wire_2), .in(wire_69), .out(wire_81));
  TC_Switch # (.UUID(64'd1362364993304987078 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_12 (.en(wire_0), .in(wire_64), .out(wire_65));
  TC_Switch # (.UUID(64'd2658338769241505139 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_13 (.en(wire_6), .in(wire_8), .out(wire_79));
  TC_Switch # (.UUID(64'd638425122573993149 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_14 (.en(wire_53), .in(wire_47), .out(wire_44));
  TC_Switch # (.UUID(64'd3619970399377026756 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_15 (.en(wire_11), .in(wire_19), .out(wire_77));
  TC_Switch # (.UUID(64'd529149196677620597 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_16 (.en(wire_32), .in(wire_19), .out(wire_36_3));
  TC_Switch # (.UUID(64'd693839758104742864 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_17 (.en(wire_17), .in(wire_47), .out(wire_36_0));
  TC_Switch # (.UUID(64'd456546521315189651 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_18 (.en(wire_29), .in(wire_8), .out(wire_36_1));
  TC_Switch # (.UUID(64'd1438168433823453622 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_19 (.en(wire_3), .in(wire_64), .out(wire_36_2));
  TC_Switch # (.UUID(64'd1745894509189344897 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_20 (.en(wire_15), .in(wire_69), .out(wire_36_4));
  TC_Switch # (.UUID(64'd916509930567616671 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_21 (.en(wire_61), .in(wire_49), .out(wire_36_5));
  TC_Switch # (.UUID(64'd2360445239048170546 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_22 (.en(wire_39), .in(wire_54), .out(wire_36_6));
  TC_Switch # (.UUID(64'd4327029652055198873 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_23 (.en(wire_9), .in(wire_20), .out(wire_36_7));
  TC_IndexerByte # (.UUID(64'd918448405620721287 ^ UUID), .INDEX(64'd0)) IndexerByte_24 (.in(wire_22), .out(wire_70));
  TC_IndexerByte # (.UUID(64'd1057721888676459279 ^ UUID), .INDEX(64'd1)) IndexerByte_25 (.in(wire_22), .out(wire_45));
  TC_IndexerByte # (.UUID(64'd1352066932906017317 ^ UUID), .INDEX(64'd2)) IndexerByte_26 (.in(wire_22), .out(wire_48));
  TC_IndexerByte # (.UUID(64'd1958548087018421884 ^ UUID), .INDEX(64'd3)) IndexerByte_27 (.in(wire_22), .out(wire_57));
  TC_IndexerByte # (.UUID(64'd1872221820076695809 ^ UUID), .INDEX(64'd4)) IndexerByte_28 (.in(wire_22), .out(wire_62));
  TC_IndexerByte # (.UUID(64'd155788635881539499 ^ UUID), .INDEX(64'd5)) IndexerByte_29 (.in(wire_22), .out(wire_59));
  TC_IndexerByte # (.UUID(64'd3607349748970436479 ^ UUID), .INDEX(64'd6)) IndexerByte_30 (.in(wire_22), .out(wire_73));
  TC_IndexerByte # (.UUID(64'd619019226309600983 ^ UUID), .INDEX(64'd7)) IndexerByte_31 (.in(wire_22), .out(wire_78));
  TC_Not # (.UUID(64'd3269442743406874800 ^ UUID), .BIT_WIDTH(64'd1)) Not_32 (.in(wire_56), .out(wire_80));
  TC_Not # (.UUID(64'd3335461814723912582 ^ UUID), .BIT_WIDTH(64'd1)) Not_33 (.in(wire_34), .out(wire_30));
  TC_Not # (.UUID(64'd2877595133194298363 ^ UUID), .BIT_WIDTH(64'd1)) Not_34 (.in(wire_63), .out(wire_74));
  TC_Not # (.UUID(64'd511029179704994023 ^ UUID), .BIT_WIDTH(64'd1)) Not_35 (.in(wire_41), .out(wire_52));
  TC_Not # (.UUID(64'd2472562442316617084 ^ UUID), .BIT_WIDTH(64'd1)) Not_36 (.in(wire_42), .out(wire_23));
  TC_Not # (.UUID(64'd2000705675645612502 ^ UUID), .BIT_WIDTH(64'd1)) Not_37 (.in(wire_31), .out(wire_37));
  TC_Not # (.UUID(64'd1452795538963522449 ^ UUID), .BIT_WIDTH(64'd1)) Not_38 (.in(wire_35), .out(wire_75));
  TC_Constant # (.UUID(64'd1586029080375720595 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_39 (.out(wire_25));
  TC_Constant # (.UUID(64'd388067972797382358 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_40 (.out(wire_55));
  TC_Constant # (.UUID(64'd1177129839986712831 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_41 (.out(wire_51));
  TC_Constant # (.UUID(64'd3356357546357843909 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_42 (.out(wire_38));
  TC_Constant # (.UUID(64'd189150637603521722 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h5)) Constant8_43 (.out(wire_60));
  TC_Constant # (.UUID(64'd325458571362803486 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_44 (.out(wire_68));
  TC_Constant # (.UUID(64'd1673740416312550615 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_45 (.out(wire_67));
  TC_Constant # (.UUID(64'd750265994278455853 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h8)) Constant8_46 (.out(wire_10));
  TC_Switch # (.UUID(64'd2313475539969607657 ^ UUID), .BIT_WIDTH(64'd64)) Output64z_47 (.en(wire_9), .in(wire_46), .out(Output));
  x10zpnz_2 # (.UUID(64'd1727933763238808163 ^ UUID)) x10zpnz_2_48 (.clk(clk), .rst(rst), .Full(wire_71), .Input(wire_40), .Output(wire_20));
  x10zpnz_2 # (.UUID(64'd2153897062672571173 ^ UUID)) x10zpnz_2_49 (.clk(clk), .rst(rst), .Full(wire_76), .Input(wire_26), .Output(wire_54));
  x10zpnz_2 # (.UUID(64'd2849872454438346445 ^ UUID)) x10zpnz_2_50 (.clk(clk), .rst(rst), .Full(wire_81), .Input(wire_72), .Output(wire_49));
  x10zpnz_2 # (.UUID(64'd2055897542852213967 ^ UUID)) x10zpnz_2_51 (.clk(clk), .rst(rst), .Full(wire_65), .Input(wire_27), .Output(wire_69));
  x10zpnz_2 # (.UUID(64'd1632279964610686668 ^ UUID)) x10zpnz_2_52 (.clk(clk), .rst(rst), .Full(wire_79), .Input(wire_4), .Output(wire_64));
  x10zpnz_2 # (.UUID(64'd3394312640399286977 ^ UUID)) x10zpnz_2_53 (.clk(clk), .rst(rst), .Full(wire_44), .Input(wire_58), .Output(wire_8));
  x10zpnz_2 # (.UUID(64'd4611331094701205989 ^ UUID)) x10zpnz_2_54 (.clk(clk), .rst(rst), .Full(wire_77), .Input(wire_18), .Output(wire_47));
  x10zpnz_2 # (.UUID(64'd1109747332268038549 ^ UUID)) x10zpnz_2_55 (.clk(clk), .rst(rst), .Full(wire_66), .Input(wire_21), .Output(wire_19));
  ByteToNumbersz_2 # (.UUID(64'd3749607521372867419 ^ UUID)) ByteToNumbersz_2_56 (.clk(clk), .rst(rst), .Input(wire_78), .Has_48(wire_14), .Number(wire_40));
  ByteToNumbersz_2 # (.UUID(64'd3913277475394169812 ^ UUID)) ByteToNumbersz_2_57 (.clk(clk), .rst(rst), .Input(wire_73), .Has_48(wire_12), .Number(wire_26));
  ByteToNumbersz_2 # (.UUID(64'd3620624112168064607 ^ UUID)) ByteToNumbersz_2_58 (.clk(clk), .rst(rst), .Input(wire_59), .Has_48(wire_7), .Number(wire_72));
  ByteToNumbersz_2 # (.UUID(64'd2323961815195874159 ^ UUID)) ByteToNumbersz_2_59 (.clk(clk), .rst(rst), .Input(wire_62), .Has_48(wire_2), .Number(wire_27));
  ByteToNumbersz_2 # (.UUID(64'd3940308161942743972 ^ UUID)) ByteToNumbersz_2_60 (.clk(clk), .rst(rst), .Input(wire_57), .Has_48(wire_0), .Number(wire_4));
  ByteToNumbersz_2 # (.UUID(64'd768896382432068357 ^ UUID)) ByteToNumbersz_2_61 (.clk(clk), .rst(rst), .Input(wire_48), .Has_48(wire_6), .Number(wire_58));
  ByteToNumbersz_2 # (.UUID(64'd3898128566190933750 ^ UUID)) ByteToNumbersz_2_62 (.clk(clk), .rst(rst), .Input(wire_45), .Has_48(wire_53), .Number(wire_18));
  ByteToNumbersz_2 # (.UUID(64'd378029805062717004 ^ UUID)) ByteToNumbersz_2_63 (.clk(clk), .rst(rst), .Input(wire_70), .Has_48(wire_11), .Number(wire_21));
  OnOrOff # (.UUID(64'd640412305280202322 ^ UUID)) OnOrOff_64 (.clk(clk), .rst(rst), .Input(wire_32), .Output(wire_56));
  OnOrOff # (.UUID(64'd4578035466279301241 ^ UUID)) OnOrOff_65 (.clk(clk), .rst(rst), .Input(wire_56), .Output(wire_34_0));
  mand # (.UUID(64'd2850811116901752460 ^ UUID)) mand_66 (.clk(clk), .rst(rst), .Input_1(wire_80), .Input_2(wire_28), .Output(wire_17));
  OnOrOff # (.UUID(64'd1212524261752792256 ^ UUID)) OnOrOff_67 (.clk(clk), .rst(rst), .Input(wire_17), .Output(wire_34_1));
  OnOrOff # (.UUID(64'd3179644437865908277 ^ UUID)) OnOrOff_68 (.clk(clk), .rst(rst), .Input(wire_34), .Output(wire_63_1));
  mand # (.UUID(64'd3277479475048403299 ^ UUID)) mand_69 (.clk(clk), .rst(rst), .Input_1(wire_30), .Input_2(wire_5), .Output(wire_29));
  OnOrOff # (.UUID(64'd2384354698056104438 ^ UUID)) OnOrOff_70 (.clk(clk), .rst(rst), .Input(wire_29), .Output(wire_63_0));
  OnOrOff # (.UUID(64'd4561424185841553039 ^ UUID)) OnOrOff_71 (.clk(clk), .rst(rst), .Input(wire_63), .Output(wire_41_0));
  mand # (.UUID(64'd4305571255693994367 ^ UUID)) mand_72 (.clk(clk), .rst(rst), .Input_1(wire_74), .Input_2(wire_13), .Output(wire_3));
  OnOrOff # (.UUID(64'd1453608781643062095 ^ UUID)) OnOrOff_73 (.clk(clk), .rst(rst), .Input(wire_3), .Output(wire_41_1));
  OnOrOff # (.UUID(64'd1582180910829622389 ^ UUID)) OnOrOff_74 (.clk(clk), .rst(rst), .Input(wire_41), .Output(wire_42_1));
  mand # (.UUID(64'd739614864554910836 ^ UUID)) mand_75 (.clk(clk), .rst(rst), .Input_1(wire_52), .Input_2(wire_24), .Output(wire_15));
  OnOrOff # (.UUID(64'd3747143776799112453 ^ UUID)) OnOrOff_76 (.clk(clk), .rst(rst), .Input(wire_15), .Output(wire_42_0));
  OnOrOff # (.UUID(64'd1280532517894966659 ^ UUID)) OnOrOff_77 (.clk(clk), .rst(rst), .Input(wire_42), .Output(wire_31_1));
  mand # (.UUID(64'd2227228807332047616 ^ UUID)) mand_78 (.clk(clk), .rst(rst), .Input_1(wire_23), .Input_2(wire_43), .Output(wire_61));
  OnOrOff # (.UUID(64'd2650310853448399114 ^ UUID)) OnOrOff_79 (.clk(clk), .rst(rst), .Input(wire_61), .Output(wire_31_0));
  OnOrOff # (.UUID(64'd1325072695741667115 ^ UUID)) OnOrOff_80 (.clk(clk), .rst(rst), .Input(wire_31), .Output(wire_35_1));
  mand # (.UUID(64'd3853908561459183764 ^ UUID)) mand_81 (.clk(clk), .rst(rst), .Input_1(wire_37), .Input_2(wire_50), .Output(wire_39));
  OnOrOff # (.UUID(64'd538149528022798750 ^ UUID)) OnOrOff_82 (.clk(clk), .rst(rst), .Input(wire_39), .Output(wire_35_0));
  OnOrOff # (.UUID(64'd2958063293918792657 ^ UUID)) OnOrOff_83 (.clk(clk), .rst(rst), .Input(wire_35), .Output(wire_33_0));
  mand # (.UUID(64'd3605908471953912169 ^ UUID)) mand_84 (.clk(clk), .rst(rst), .Input_1(wire_75), .Input_2(wire_16), .Output(wire_9));
  OnOrOff # (.UUID(64'd4050520338198485190 ^ UUID)) OnOrOff_85 (.clk(clk), .rst(rst), .Input(wire_9), .Output(wire_33_1));
  _8rSwitch # (.UUID(64'd3759739111363517803 ^ UUID)) _8rSwitch_86 (.clk(clk), .rst(rst), .Enable(wire_32), .Input(wire_25), .Output(wire_1_7));
  _8rSwitch # (.UUID(64'd3050627992690140294 ^ UUID)) _8rSwitch_87 (.clk(clk), .rst(rst), .Enable(wire_17), .Input(wire_55), .Output(wire_1_6));
  _8rSwitch # (.UUID(64'd4012340497973258837 ^ UUID)) _8rSwitch_88 (.clk(clk), .rst(rst), .Enable(wire_29), .Input(wire_51), .Output(wire_1_5));
  _8rSwitch # (.UUID(64'd2776943117159413848 ^ UUID)) _8rSwitch_89 (.clk(clk), .rst(rst), .Enable(wire_3), .Input(wire_38), .Output(wire_1_4));
  _8rSwitch # (.UUID(64'd2151440494668335396 ^ UUID)) _8rSwitch_90 (.clk(clk), .rst(rst), .Enable(wire_15), .Input(wire_60), .Output(wire_1_3));
  _8rSwitch # (.UUID(64'd2638808000486651592 ^ UUID)) _8rSwitch_91 (.clk(clk), .rst(rst), .Enable(wire_61), .Input(wire_68), .Output(wire_1_2));
  _8rSwitch # (.UUID(64'd1123854421980830513 ^ UUID)) _8rSwitch_92 (.clk(clk), .rst(rst), .Enable(wire_39), .Input(wire_67), .Output(wire_1_1));
  _8rSwitch # (.UUID(64'd1020953886359072499 ^ UUID)) _8rSwitch_93 (.clk(clk), .rst(rst), .Enable(wire_9), .Input(wire_10), .Output(wire_1_0));

  wire [0:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_1_0;
  wire [7:0] wire_1_1;
  wire [7:0] wire_1_2;
  wire [7:0] wire_1_3;
  wire [7:0] wire_1_4;
  wire [7:0] wire_1_5;
  wire [7:0] wire_1_6;
  wire [7:0] wire_1_7;
  assign wire_1 = wire_1_0|wire_1_1|wire_1_2|wire_1_3|wire_1_4|wire_1_5|wire_1_6|wire_1_7;
  assign Offset = wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [63:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [7:0] wire_18;
  wire [63:0] wire_19;
  wire [63:0] wire_20;
  wire [7:0] wire_21;
  wire [63:0] wire_22;
  assign wire_22 = Main_8b;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [7:0] wire_25;
  wire [7:0] wire_26;
  wire [7:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_31_0;
  wire [0:0] wire_31_1;
  assign wire_31 = wire_31_0|wire_31_1;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_33_0;
  wire [0:0] wire_33_1;
  assign wire_33 = wire_33_0|wire_33_1;
  wire [0:0] wire_34;
  wire [0:0] wire_34_0;
  wire [0:0] wire_34_1;
  assign wire_34 = wire_34_0|wire_34_1;
  wire [0:0] wire_35;
  wire [0:0] wire_35_0;
  wire [0:0] wire_35_1;
  assign wire_35 = wire_35_0|wire_35_1;
  wire [63:0] wire_36;
  wire [63:0] wire_36_0;
  wire [63:0] wire_36_1;
  wire [63:0] wire_36_2;
  wire [63:0] wire_36_3;
  wire [63:0] wire_36_4;
  wire [63:0] wire_36_5;
  wire [63:0] wire_36_6;
  wire [63:0] wire_36_7;
  assign wire_36 = wire_36_0|wire_36_1|wire_36_2|wire_36_3|wire_36_4|wire_36_5|wire_36_6|wire_36_7;
  assign Value = wire_36;
  wire [0:0] wire_37;
  wire [7:0] wire_38;
  wire [0:0] wire_39;
  wire [7:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_41_0;
  wire [0:0] wire_41_1;
  assign wire_41 = wire_41_0|wire_41_1;
  wire [0:0] wire_42;
  wire [0:0] wire_42_0;
  wire [0:0] wire_42_1;
  assign wire_42 = wire_42_0|wire_42_1;
  wire [0:0] wire_43;
  wire [63:0] wire_44;
  wire [7:0] wire_45;
  wire [63:0] wire_46;
  wire [63:0] wire_47;
  wire [7:0] wire_48;
  wire [63:0] wire_49;
  wire [0:0] wire_50;
  wire [7:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [63:0] wire_54;
  wire [7:0] wire_55;
  wire [0:0] wire_56;
  wire [7:0] wire_57;
  wire [7:0] wire_58;
  wire [7:0] wire_59;
  wire [7:0] wire_60;
  wire [0:0] wire_61;
  wire [7:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_63_0;
  wire [0:0] wire_63_1;
  assign wire_63 = wire_63_0|wire_63_1;
  wire [63:0] wire_64;
  wire [63:0] wire_65;
  wire [63:0] wire_66;
  assign wire_66 = Carry_In;
  wire [7:0] wire_67;
  wire [7:0] wire_68;
  wire [63:0] wire_69;
  wire [7:0] wire_70;
  wire [63:0] wire_71;
  wire [7:0] wire_72;
  wire [7:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [63:0] wire_76;
  wire [63:0] wire_77;
  wire [7:0] wire_78;
  wire [63:0] wire_79;
  wire [0:0] wire_80;
  wire [63:0] wire_81;

endmodule
