module is0 (clk, rst, Input, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [15:0] Input;
  output  wire [0:0] Output;

  TC_Splitter16 # (.UUID(64'd2172339877071428244 ^ UUID)) Splitter16_0 (.in(wire_6), .out0(wire_17), .out1(wire_12));
  TC_Splitter8 # (.UUID(64'd4068030003329438922 ^ UUID)) Splitter8_1 (.in(wire_12), .out0(wire_4), .out1(wire_7), .out2(wire_15), .out3(wire_9), .out4(wire_19), .out5(wire_16), .out6(wire_14), .out7(wire_2));
  TC_Splitter8 # (.UUID(64'd4301914091385864416 ^ UUID)) Splitter8_2 (.in(wire_17), .out0(wire_5), .out1(wire_8), .out2(wire_18), .out3(wire_10), .out4(wire_20), .out5(wire_13), .out6(wire_11), .out7(wire_3));
  OnOrOff # (.UUID(64'd2324880171805938053 ^ UUID)) OnOrOff_3 (.clk(clk), .rst(rst), .Input(wire_5), .Output(wire_1_15));
  OnOrOff # (.UUID(64'd888330152005551935 ^ UUID)) OnOrOff_4 (.clk(clk), .rst(rst), .Input(wire_8), .Output(wire_1_14));
  OnOrOff # (.UUID(64'd2336601701524891901 ^ UUID)) OnOrOff_5 (.clk(clk), .rst(rst), .Input(wire_18), .Output(wire_1_13));
  OnOrOff # (.UUID(64'd3144173771624457841 ^ UUID)) OnOrOff_6 (.clk(clk), .rst(rst), .Input(wire_10), .Output(wire_1_12));
  OnOrOff # (.UUID(64'd2211053769255465488 ^ UUID)) OnOrOff_7 (.clk(clk), .rst(rst), .Input(wire_20), .Output(wire_1_11));
  OnOrOff # (.UUID(64'd4188011463506493338 ^ UUID)) OnOrOff_8 (.clk(clk), .rst(rst), .Input(wire_13), .Output(wire_1_9));
  OnOrOff # (.UUID(64'd3485928475127179510 ^ UUID)) OnOrOff_9 (.clk(clk), .rst(rst), .Input(wire_3), .Output(wire_1_5));
  OnOrOff # (.UUID(64'd1049174922350773654 ^ UUID)) OnOrOff_10 (.clk(clk), .rst(rst), .Input(wire_11), .Output(wire_1_7));
  OnOrOff # (.UUID(64'd4441576353850611950 ^ UUID)) OnOrOff_11 (.clk(clk), .rst(rst), .Input(wire_4), .Output(wire_1_3));
  OnOrOff # (.UUID(64'd4487118609378894987 ^ UUID)) OnOrOff_12 (.clk(clk), .rst(rst), .Input(wire_7), .Output(wire_1_0));
  OnOrOff # (.UUID(64'd3315847775754123915 ^ UUID)) OnOrOff_13 (.clk(clk), .rst(rst), .Input(wire_15), .Output(wire_1_1));
  OnOrOff # (.UUID(64'd2288588140048734080 ^ UUID)) OnOrOff_14 (.clk(clk), .rst(rst), .Input(wire_19), .Output(wire_1_4));
  OnOrOff # (.UUID(64'd2792623782746976428 ^ UUID)) OnOrOff_15 (.clk(clk), .rst(rst), .Input(wire_2), .Output(wire_1_10));
  OnOrOff # (.UUID(64'd3437272793363400400 ^ UUID)) OnOrOff_16 (.clk(clk), .rst(rst), .Input(wire_14), .Output(wire_1_8));
  OnOrOff # (.UUID(64'd1820009483342798816 ^ UUID)) OnOrOff_17 (.clk(clk), .rst(rst), .Input(wire_16), .Output(wire_1_6));
  OnOrOff # (.UUID(64'd3062162042557451159 ^ UUID)) OnOrOff_18 (.clk(clk), .rst(rst), .Input(wire_9), .Output(wire_1_2));
  TC_Not # (.UUID(64'd573715845666441797 ^ UUID), .BIT_WIDTH(64'd1)) Not_19 (.in(wire_1), .out(wire_0));

  wire [0:0] wire_0;
  assign Output = wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_1_0;
  wire [0:0] wire_1_1;
  wire [0:0] wire_1_2;
  wire [0:0] wire_1_3;
  wire [0:0] wire_1_4;
  wire [0:0] wire_1_5;
  wire [0:0] wire_1_6;
  wire [0:0] wire_1_7;
  wire [0:0] wire_1_8;
  wire [0:0] wire_1_9;
  wire [0:0] wire_1_10;
  wire [0:0] wire_1_11;
  wire [0:0] wire_1_12;
  wire [0:0] wire_1_13;
  wire [0:0] wire_1_14;
  wire [0:0] wire_1_15;
  assign wire_1 = wire_1_0|wire_1_1|wire_1_2|wire_1_3|wire_1_4|wire_1_5|wire_1_6|wire_1_7|wire_1_8|wire_1_9|wire_1_10|wire_1_11|wire_1_12|wire_1_13|wire_1_14|wire_1_15;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [15:0] wire_6;
  assign wire_6 = Input;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [7:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [7:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;

endmodule
