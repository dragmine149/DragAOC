module RangeChecker (clk, rst, Input_1, Input_2, Input_3, Input_4, Input_5, Input_6, Input_7, Input_8, Input_9, Input_10, Input_11, Input_12, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Input_1;
  input  wire [7:0] Input_2;
  input  wire [7:0] Input_3;
  input  wire [7:0] Input_4;
  input  wire [7:0] Input_5;
  input  wire [7:0] Input_6;
  input  wire [7:0] Input_7;
  input  wire [7:0] Input_8;
  input  wire [7:0] Input_9;
  input  wire [7:0] Input_10;
  input  wire [7:0] Input_11;
  input  wire [7:0] Input_12;
  output  wire [0:0] Output;

  TC_LessI # (.UUID(64'd17102259344944258 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_0 (.in0(wire_15), .in1(wire_7), .out(wire_19));
  TC_Equal # (.UUID(64'd2880193297870243694 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_1 (.in0(wire_15), .in1(wire_7), .out(wire_21));
  TC_Switch # (.UUID(64'd2429876860692029960 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_2 (.en(wire_19), .in(wire_19), .out(wire_4_4));
  TC_LessI # (.UUID(64'd3237086543786144998 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_3 (.in0(wire_20), .in1(wire_2), .out(wire_29));
  TC_Equal # (.UUID(64'd2333243112151950960 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_4 (.in0(wire_20), .in1(wire_2), .out(wire_27));
  TC_And # (.UUID(64'd495205846149705491 ^ UUID), .BIT_WIDTH(64'd1)) And_5 (.in0(wire_21), .in1(wire_29), .out(wire_5));
  TC_Switch # (.UUID(64'd1852381923696279992 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_6 (.en(wire_5), .in(wire_5), .out(wire_4_5));
  TC_LessI # (.UUID(64'd1396085881594691849 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_7 (.in0(wire_0), .in1(wire_3), .out(wire_22));
  TC_Equal # (.UUID(64'd1412372811851921160 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_8 (.in0(wire_0), .in1(wire_3), .out(wire_28));
  TC_And # (.UUID(64'd439381512683118739 ^ UUID), .BIT_WIDTH(64'd1)) And_9 (.in0(wire_25), .in1(wire_22), .out(wire_18));
  TC_Switch # (.UUID(64'd2119929393328876927 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_10 (.en(wire_18), .in(wire_18), .out(wire_4_3));
  TC_LessI # (.UUID(64'd1342297543562718294 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_11 (.in0(wire_12), .in1(wire_17), .out(wire_10));
  TC_Equal # (.UUID(64'd2466326283072686500 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_12 (.in0(wire_12), .in1(wire_17), .out(wire_32));
  TC_And # (.UUID(64'd1821600307067016021 ^ UUID), .BIT_WIDTH(64'd1)) And_13 (.in0(wire_1), .in1(wire_10), .out(wire_14));
  TC_Switch # (.UUID(64'd2029728654402094425 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_14 (.en(wire_14), .in(wire_14), .out(wire_4_2));
  TC_LessI # (.UUID(64'd2661190807025871762 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_15 (.in0(wire_26), .in1(wire_11), .out(wire_6));
  TC_Equal # (.UUID(64'd605369283700856452 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_16 (.in0(wire_26), .in1(wire_11), .out(wire_24));
  TC_And # (.UUID(64'd814807313563712626 ^ UUID), .BIT_WIDTH(64'd1)) And_17 (.in0(wire_31), .in1(wire_6), .out(wire_13));
  TC_Switch # (.UUID(64'd3597646569637874046 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_18 (.en(wire_13), .in(wire_13), .out(wire_4_0));
  TC_LessI # (.UUID(64'd2893908673290003885 ^ UUID), .BIT_WIDTH(64'd8)) LessI8_19 (.in0(wire_16), .in1(wire_9), .out(wire_23));
  TC_Equal # (.UUID(64'd3417917873528509733 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_20 (.in0(wire_16), .in1(wire_9), .out());
  TC_And # (.UUID(64'd262212562981118540 ^ UUID), .BIT_WIDTH(64'd1)) And_21 (.in0(wire_30), .in1(wire_23), .out(wire_8));
  TC_Switch # (.UUID(64'd1928959780033807708 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_22 (.en(wire_8), .in(wire_8), .out(wire_4_1));
  TC_Constant # (.UUID(64'd3882103631809293241 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_23 (.out());
  TC_Constant # (.UUID(64'd433799539696246386 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_24 (.out());
  TC_Constant # (.UUID(64'd2026647646301893397 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_25 (.out());
  TC_Constant # (.UUID(64'd3007645625930056830 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_26 (.out());
  TC_Constant # (.UUID(64'd3680454433287952494 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_27 (.out());
  TC_Switch # (.UUID(64'd3023000740973880929 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_28 (.en(wire_5), .in(wire_27), .out(wire_25));
  TC_Switch # (.UUID(64'd3127937551302518160 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_29 (.en(wire_18), .in(wire_28), .out(wire_1));
  TC_Switch # (.UUID(64'd2978497890833559325 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_30 (.en(wire_14), .in(wire_32), .out(wire_31));
  TC_Switch # (.UUID(64'd4241732967994556158 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_31 (.en(wire_13), .in(wire_24), .out(wire_30));

  wire [7:0] wire_0;
  assign wire_0 = Input_11;
  wire [0:0] wire_1;
  wire [7:0] wire_2;
  assign wire_2 = Input_2;
  wire [7:0] wire_3;
  assign wire_3 = Input_12;
  wire [0:0] wire_4;
  wire [0:0] wire_4_0;
  wire [0:0] wire_4_1;
  wire [0:0] wire_4_2;
  wire [0:0] wire_4_3;
  wire [0:0] wire_4_4;
  wire [0:0] wire_4_5;
  assign wire_4 = wire_4_0|wire_4_1|wire_4_2|wire_4_3|wire_4_4|wire_4_5;
  assign Output = wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [7:0] wire_7;
  assign wire_7 = Input_4;
  wire [0:0] wire_8;
  wire [7:0] wire_9;
  assign wire_9 = Input_6;
  wire [0:0] wire_10;
  wire [7:0] wire_11;
  assign wire_11 = Input_8;
  wire [7:0] wire_12;
  assign wire_12 = Input_9;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [7:0] wire_15;
  assign wire_15 = Input_3;
  wire [7:0] wire_16;
  assign wire_16 = Input_5;
  wire [7:0] wire_17;
  assign wire_17 = Input_10;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [7:0] wire_20;
  assign wire_20 = Input_1;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [7:0] wire_26;
  assign wire_26 = Input_7;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;

endmodule
