module Day2Part2 (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_Constant # (.UUID(64'd1726993617052590723 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFFFFFFFFFFFFFFFF)) Constant64_0 (.out(wire_101));
  TC_FileLoader # (.UUID(64'd3987767967543158583 ^ UUID), .DEFAULT_FILE_NAME("day2_modified")) FileLoader_1 (.clk(clk), .rst(rst), .en(wire_32), .address(wire_0), .out(wire_35_0));
  TC_Constant # (.UUID(64'd337803116546834142 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_2 (.out(wire_32));
  TC_LessU # (.UUID(64'd2415299641673726094 ^ UUID), .BIT_WIDTH(64'd64)) LessU64_3 (.in0(wire_59), .in1(wire_0), .out(wire_37));
  TC_FileLoader # (.UUID(64'd4235385288069024156 ^ UUID), .DEFAULT_FILE_NAME("day2_test_1")) FileLoader_4 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_0), .out(wire_35_1));
  TC_Constant # (.UUID(64'd1484234401691717814 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_5 (.out());
  TC_DelayLine # (.UUID(64'd2141883989358176841 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_6 (.clk(clk), .rst(rst), .in(wire_12), .out(wire_90));
  TC_Add # (.UUID(64'd3665390526026043059 ^ UUID), .BIT_WIDTH(64'd64)) Add64_7 (.in0({{56{1'b0}}, wire_6 }), .in1(wire_0), .ci(1'd0), .out(wire_57), .co());
  TC_Counter # (.UUID(64'd3781882184507484018 ^ UUID), .BIT_WIDTH(64'd64), .count(64'd1)) Counter64_8 (.clk(clk), .rst(rst), .save(wire_83), .in(wire_14), .out(wire_5));
  TC_Not # (.UUID(64'd2915069602117248147 ^ UUID), .BIT_WIDTH(64'd1)) Not_9 (.in(wire_37), .out(wire_25));
  TC_And # (.UUID(64'd4444366698480428793 ^ UUID), .BIT_WIDTH(64'd1)) And_10 (.in0(wire_61), .in1(wire_37), .out(wire_42));
  TC_Or # (.UUID(64'd1455535717111312185 ^ UUID), .BIT_WIDTH(64'd1)) Or_11 (.in0(wire_34), .in1(wire_42), .out(wire_83));
  TC_Not # (.UUID(64'd4292279915901693506 ^ UUID), .BIT_WIDTH(64'd1)) Not_12 (.in(wire_61), .out(wire_34));
  TC_Switch # (.UUID(64'd259253643073170517 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_13 (.en(wire_25), .in(wire_5), .out(wire_19_1));
  TC_Counter # (.UUID(64'd4027361701724138616 ^ UUID), .BIT_WIDTH(64'd64), .count(64'd1)) Counter64_14 (.clk(clk), .rst(rst), .save(wire_78), .in(wire_58), .out(wire_44));
  TC_Ram # (.UUID(64'd3231836939472590219 ^ UUID), .WORD_WIDTH(64'd64), .WORD_COUNT(64'd1250)) Ram_15 (.clk(clk), .rst(rst), .load(wire_89), .save(wire_40), .address(wire_9[31:0]), .in0(wire_98), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_18), .out1(), .out2(), .out3());
  TC_Halt # (.UUID(64'd1646709671390234641 ^ UUID), .HALT_MESSAGE("Program finished!")) Halt_16 (.clk(clk), .rst(rst), .en(wire_72));
  TC_NoteSound # (.UUID(64'd2856162216424263791 ^ UUID)) NoteSound_17 (.clk(clk), .rst(rst), .command({{7{1'b0}}, wire_72 }), .note(wire_54), .pitch(8'd0));
  TC_Constant # (.UUID(64'd3448097267265053438 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h28)) Constant8_18 (.out(wire_54));
  TC_Not # (.UUID(64'd1023328388184503186 ^ UUID), .BIT_WIDTH(64'd1)) Not_19 (.in(wire_42), .out(wire_104));
  TC_DelayLine # (.UUID(64'd4092965687359902133 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_20 (.clk(clk), .rst(rst), .in(wire_70), .out(wire_49));
  TC_Mux # (.UUID(64'd316725708318265243 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_21 (.sel(wire_61), .in0(wire_101), .in1(wire_49), .out(wire_0));
  TC_Switch # (.UUID(64'd3903258603175327041 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_22 (.en(wire_1), .in(wire_18), .out(wire_22));
  TC_Switch # (.UUID(64'd1710097796709442780 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_23 (.en(wire_8), .in(wire_18), .out(wire_30));
  TC_Switch # (.UUID(64'd3052143593441878759 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_24 (.en(wire_38), .in(wire_47), .out(wire_19_3));
  TC_Constant # (.UUID(64'd3240501465042579115 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_25 (.out(wire_87));
  TC_Not # (.UUID(64'd1867582932362601439 ^ UUID), .BIT_WIDTH(64'd1)) Not_26 (.in(wire_78), .out(wire_53));
  TC_DelayLine # (.UUID(64'd2677504830674658084 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_27 (.clk(clk), .rst(rst), .in(wire_93), .out(wire_66));
  TC_Switch # (.UUID(64'd1725179244806057793 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_28 (.en(wire_76), .in(wire_22), .out(wire_93));
  TC_DelayLine # (.UUID(64'd1784992797701007900 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_29 (.clk(clk), .rst(rst), .in(wire_76), .out(wire_55));
  TC_DelayLine # (.UUID(64'd4350311000933170162 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_30 (.clk(clk), .rst(rst), .in(wire_8), .out(wire_15));
  TC_Switch # (.UUID(64'd4182440545682965520 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_31 (.en(wire_46), .in(wire_30), .out(wire_56));
  TC_DelayLine # (.UUID(64'd247377800554737393 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_32 (.clk(clk), .rst(rst), .in(wire_56), .out(wire_41));
  TC_DelayLine # (.UUID(64'd3700638478856170501 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_33 (.clk(clk), .rst(rst), .in(wire_46), .out(wire_92));
  TC_Switch # (.UUID(64'd3804153078929315197 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_34 (.en(wire_55), .in(wire_66), .out(wire_47_1));
  TC_Switch # (.UUID(64'd79719301686403854 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_35 (.en(wire_92), .in(wire_41), .out(wire_47_0));
  TC_Add # (.UUID(64'd1069550484725226130 ^ UUID), .BIT_WIDTH(64'd64)) Add64_36 (.in0(wire_43), .in1(wire_16), .ci(1'd0), .out(wire_77), .co());
  TC_Mul # (.UUID(64'd924182476717345043 ^ UUID), .BIT_WIDTH(64'd64)) Mul64_37 (.in0(wire_43), .in1(wire_16), .out0(wire_33), .out1());
  TC_Switch # (.UUID(64'd935510424511562668 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_38 (.en(wire_75), .in(wire_77), .out(wire_67_1));
  TC_Switch # (.UUID(64'd3389748284807452395 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_39 (.en(wire_21), .in(wire_33), .out(wire_67_0));
  TC_Halt # (.UUID(64'd3795677300099293191 ^ UUID), .HALT_MESSAGE("Opcode 99 Reached!")) Halt_40 (.clk(clk), .rst(rst), .en(1'd0));
  TC_Switch # (.UUID(64'd1224855048361981157 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_41 (.en(wire_17), .in(wire_67), .out(wire_4_1));
  TC_And # (.UUID(64'd4423175184107256786 ^ UUID), .BIT_WIDTH(64'd1)) And_42 (.in0(wire_73), .in1(wire_3), .out(wire_17));
  TC_Constant # (.UUID(64'd2201783711648500038 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_43 (.out(wire_3));
  TC_Not # (.UUID(64'd3940936562307563579 ^ UUID), .BIT_WIDTH(64'd1)) Not_44 (.in(wire_17), .out(wire_102));
  TC_DelayLine # (.UUID(64'd366563469061908473 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_45 (.clk(clk), .rst(rst), .in(wire_102), .out(wire_108));
  TC_Not # (.UUID(64'd23546066323564917 ^ UUID), .BIT_WIDTH(64'd1)) Not_46 (.in(wire_42), .out(wire_95));
  TC_Or3 # (.UUID(64'd1565632499214780517 ^ UUID), .BIT_WIDTH(64'd1)) Or3_47 (.in0(wire_38), .in1(wire_79), .in2(wire_104), .out(wire_78_1));
  TC_Not # (.UUID(64'd601742535760828746 ^ UUID), .BIT_WIDTH(64'd1)) Not_48 (.in(wire_109), .out(wire_10));
  TC_DelayLine # (.UUID(64'd1263282884327671549 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_49 (.clk(clk), .rst(rst), .in(wire_1), .out(wire_26));
  TC_Not # (.UUID(64'd4567426784455268513 ^ UUID), .BIT_WIDTH(64'd1)) Not_50 (.in(wire_26), .out(wire_31));
  TC_Not # (.UUID(64'd4522425577002129070 ^ UUID), .BIT_WIDTH(64'd1)) Not_51 (.in(wire_15), .out(wire_96));
  TC_Or # (.UUID(64'd571059853550174113 ^ UUID), .BIT_WIDTH(64'd1)) Or_52 (.in0(wire_20), .in1(wire_17), .out(wire_79));
  TC_FileLoader # (.UUID(64'd4032583951989155851 ^ UUID), .DEFAULT_FILE_NAME("day2_test_2")) FileLoader_53 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_0), .out(wire_35_2));
  TC_Constant # (.UUID(64'd1883781277529937826 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_54 (.out());
  TC_Constant # (.UUID(64'd4566527038733230091 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_55 (.out());
  TC_Constant # (.UUID(64'd3138890809031518109 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_56 (.out());
  TC_Constant # (.UUID(64'd2829021048917779791 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_57 (.out());
  TC_Constant # (.UUID(64'd1405985673201260239 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_58 (.out());
  TC_Constant # (.UUID(64'd3716163551666950261 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_59 (.out());
  TC_Constant # (.UUID(64'd4023943151529497828 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_60 (.out());
  TC_Constant # (.UUID(64'd2532988701438288488 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_61 (.out());
  TC_Constant # (.UUID(64'd4214058095318520776 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_62 (.out());
  TC_Constant # (.UUID(64'd958940107339709111 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_63 (.out());
  TC_Constant # (.UUID(64'd2113422115012713154 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_64 (.out());
  TC_Constant # (.UUID(64'd372203303927728035 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_65 (.out());
  TC_Constant # (.UUID(64'd4215445727210423365 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_66 (.out());
  TC_Constant # (.UUID(64'd4177145269316879433 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_67 (.out());
  TC_FileLoader # (.UUID(64'd3305349617174586722 ^ UUID), .DEFAULT_FILE_NAME("day2_test_3")) FileLoader_68 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_0), .out(wire_35_3));
  TC_FileLoader # (.UUID(64'd231382507668522051 ^ UUID), .DEFAULT_FILE_NAME("day2_test_4")) FileLoader_69 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_0), .out(wire_35_4));
  TC_FileLoader # (.UUID(64'd1231532553883646540 ^ UUID), .DEFAULT_FILE_NAME("day2_test_5")) FileLoader_70 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_0), .out(wire_35_5));
  TC_Equal # (.UUID(64'd2821604189245118802 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_71 (.in0(wire_5), .in1({{56{1'b0}}, wire_110 }), .out(wire_52));
  TC_Equal # (.UUID(64'd834176164977634459 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_72 (.in0(wire_5), .in1({{56{1'b0}}, wire_99 }), .out(wire_86));
  TC_Constant # (.UUID(64'd1065572658605867570 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_73 (.out(wire_110));
  TC_Constant # (.UUID(64'd991865579609327770 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_74 (.out(wire_99));
  TC_Switch # (.UUID(64'd1746571703522486786 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_75 (.en(wire_52), .in(wire_80), .out(wire_23_0));
  TC_Switch # (.UUID(64'd1454525939490593477 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_76 (.en(wire_86), .in(wire_88), .out(wire_23_1));
  TC_Switch # (.UUID(64'd1728873000476622687 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_77 (.en(wire_68), .in(wire_94[7:0]), .out(wire_23_2));
  TC_Nor # (.UUID(64'd4535549015773012659 ^ UUID), .BIT_WIDTH(64'd1)) Nor_78 (.in0(wire_52), .in1(wire_86), .out(wire_68));
  TC_Equal # (.UUID(64'd4382296156982196310 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_79 (.in0(wire_18), .in1(wire_82), .out(wire_85));
  TC_And # (.UUID(64'd1888702582889417503 ^ UUID), .BIT_WIDTH(64'd1)) And_80 (.in0(wire_85), .in1(wire_20), .out(wire_65));
  TC_Halt # (.UUID(64'd4563628704689697466 ^ UUID), .HALT_MESSAGE("Number pair found!")) Halt_81 (.clk(clk), .rst(rst), .en(wire_65));
  TC_Constant # (.UUID(64'd2825119468061589370 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h12C74E0)) Constant64_82 (.out(wire_82));
  TC_Counter # (.UUID(64'd3716028370518343304 ^ UUID), .BIT_WIDTH(64'd64), .count(64'd1)) Counter64_83 (.clk(clk), .rst(rst), .save(wire_28), .in(64'd0), .out(wire_51));
  TC_Equal # (.UUID(64'd1232986498560230343 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_84 (.in0(wire_51), .in1(wire_5), .out(wire_45));
  TC_Not # (.UUID(64'd636674039187011040 ^ UUID), .BIT_WIDTH(64'd1)) Not_85 (.in(wire_7), .out(wire_28));
  TC_And # (.UUID(64'd2718161313928938546 ^ UUID), .BIT_WIDTH(64'd1)) And_86 (.in0(wire_7), .in1(wire_11), .out(wire_62));
  TC_Switch # (.UUID(64'd881720095141849915 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_87 (.en(wire_62), .in(wire_51), .out(wire_9_1));
  TC_Not # (.UUID(64'd913028056677067501 ^ UUID), .BIT_WIDTH(64'd1)) Not_88 (.in(wire_62), .out(wire_13));
  TC_Not # (.UUID(64'd952276765596778979 ^ UUID), .BIT_WIDTH(64'd1)) Not_89 (.in(wire_45), .out(wire_11));
  TC_Switch # (.UUID(64'd2786939255044915453 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_90 (.en(wire_24), .in(wire_5), .out(wire_14));
  TC_DelayLine # (.UUID(64'd333550580747512898 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_91 (.clk(clk), .rst(rst), .in(wire_62), .out(wire_81));
  TC_Halt # (.UUID(64'd173880931492206516 ^ UUID), .HALT_MESSAGE("Memory Cleared")) Halt_92 (.clk(clk), .rst(rst), .en(1'd0));
  TC_And # (.UUID(64'd1254581417745991036 ^ UUID), .BIT_WIDTH(64'd1)) And_93 (.in0(wire_48), .in1(wire_45), .out(wire_27));
  TC_Switch # (.UUID(64'd2236419431862390674 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_94 (.en(wire_24), .in(wire_57), .out(wire_70));
  TC_Not # (.UUID(64'd895591967131792673 ^ UUID), .BIT_WIDTH(64'd1)) Not_95 (.in(wire_27), .out(wire_24));
  TC_Switch # (.UUID(64'd1341671548569791167 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_96 (.en(wire_39), .in(wire_44), .out(wire_58));
  TC_DelayLine # (.UUID(64'd71778258165389772 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_97 (.clk(clk), .rst(rst), .in(wire_20), .out(wire_100));
  TC_Not # (.UUID(64'd1026398734405901705 ^ UUID), .BIT_WIDTH(64'd1)) Not_98 (.in(wire_39), .out(wire_91));
  TC_DelayLine # (.UUID(64'd3662433804087744831 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_99 (.clk(clk), .rst(rst), .in(wire_24), .out(wire_39));
  TC_Halt # (.UUID(64'd2336335384836364761 ^ UUID), .HALT_MESSAGE("Panic! Not found number within time frame!")) Halt_100 (.clk(clk), .rst(rst), .en(wire_106));
  QuickSave # (.UUID(64'd2695330121804011308 ^ UUID)) QuickSave_101 (.clk(clk), .rst(rst), .Value(wire_35), .\Number_(stored) (wire_59), .\Saved?_1 (wire_61), .\Saved?_2 ());
  BytesToNumbersz_3 # (.UUID(64'd1729469431074511873 ^ UUID)) BytesToNumbersz_3_102 (.clk(clk), .rst(rst), .Main_8b(wire_35), .Carry_In(wire_90), .Output(wire_12), .Offset(wire_6), .Value(wire_94));
  OnOrOff # (.UUID(64'd3163142382288365090 ^ UUID)) OnOrOff_103 (.clk(clk), .rst(rst), .Input(wire_25), .Output(wire_2_1));
  flippedzm64bzmswitch # (.UUID(64'd2031059029553199162 ^ UUID)) flippedzm64bzmswitch_104 (.clk(clk), .rst(rst), .Input_1(wire_44), .Input_2(wire_53), .Output(wire_19_0));
  OnOrOff # (.UUID(64'd150349705086353648 ^ UUID)) OnOrOff_105 (.clk(clk), .rst(rst), .Input(wire_53), .Output(wire_29_1));
  OnOrOff # (.UUID(64'd224193335304047014 ^ UUID)) OnOrOff_106 (.clk(clk), .rst(rst), .Input(wire_103), .Output(wire_29_2));
  mand # (.UUID(64'd3349436745291189726 ^ UUID)) mand_107 (.clk(clk), .rst(rst), .Input_1(wire_38), .Input_2(wire_87), .Output(wire_103));
  mand # (.UUID(64'd242248694494001734 ^ UUID)) mand_108 (.clk(clk), .rst(rst), .Input_1(wire_42), .Input_2(wire_108), .Output(wire_109));
  flippedzm64bzmswitch # (.UUID(64'd1881707450118815654 ^ UUID)) flippedzm64bzmswitch_109 (.clk(clk), .rst(rst), .Input_1(wire_22), .Input_2(wire_26), .Output(wire_71));
  OnOrOff # (.UUID(64'd4158355321388927517 ^ UUID)) OnOrOff_110 (.clk(clk), .rst(rst), .Input(wire_55), .Output(wire_38_0));
  flippedzm64bzmswitch # (.UUID(64'd558922318308219109 ^ UUID)) flippedzm64bzmswitch_111 (.clk(clk), .rst(rst), .Input_1(wire_30), .Input_2(wire_15), .Output(wire_63));
  OnOrOff # (.UUID(64'd3868852299644989347 ^ UUID)) OnOrOff_112 (.clk(clk), .rst(rst), .Input(wire_92), .Output(wire_38_1));
  Opcodez_zmz_1z_2z_99 # (.UUID(64'd1253066027045582023 ^ UUID)) Opcodez_zmz_1z_2z_99_113 (.clk(clk), .rst(rst), .Opcode(wire_69[7:0]), .Add(wire_75), .divide(wire_21), .halt(wire_20));
  OnOrOff # (.UUID(64'd779081389060044986 ^ UUID)) OnOrOff_114 (.clk(clk), .rst(rst), .Input(wire_17), .Output(wire_2_0));
  flippedzm64bzmswitch # (.UUID(64'd3330710435434371616 ^ UUID)) flippedzm64bzmswitch_115 (.clk(clk), .rst(rst), .Input_1(wire_60), .Input_2(wire_17), .Output(wire_19_2));
  flippedzm64bzmswitch # (.UUID(64'd3395453474976780481 ^ UUID)) flippedzm64bzmswitch_116 (.clk(clk), .rst(rst), .Input_1({{56{1'b0}}, wire_23 }), .Input_2(wire_95), .Output(wire_4_0));
  CellWritter # (.UUID(64'd1760994904368207804 ^ UUID)) CellWritter_117 (.clk(clk), .rst(rst), .Clear(wire_10), .Write(wire_29), .Value_1(wire_18), .Value_2(wire_69), .Written(wire_97));
  CellWritter # (.UUID(64'd2225673571882546958 ^ UUID)) CellWritter_118 (.clk(clk), .rst(rst), .Clear(wire_10), .Write(wire_26), .Value_1(wire_71), .Value_2(wire_43), .Written(wire_64));
  CellWritter # (.UUID(64'd640733034693975124 ^ UUID)) CellWritter_119 (.clk(clk), .rst(rst), .Clear(wire_10), .Write(wire_15), .Value_1(wire_63), .Value_2(wire_16), .Written(wire_50));
  mand # (.UUID(64'd2253745888330672149 ^ UUID)) mand_120 (.clk(clk), .rst(rst), .Input_1(wire_1), .Input_2(wire_31), .Output(wire_76));
  mand # (.UUID(64'd4089700112481536660 ^ UUID)) mand_121 (.clk(clk), .rst(rst), .Input_1(wire_8), .Input_2(wire_96), .Output(wire_46));
  CellWritter # (.UUID(64'd3735606448599014512 ^ UUID)) CellWritter_122 (.clk(clk), .rst(rst), .Clear(wire_10), .Write(wire_74), .Value_1(wire_18), .Value_2(wire_60), .Written(wire_73));
  mand # (.UUID(64'd1207172339067544539 ^ UUID)) mand_123 (.clk(clk), .rst(rst), .Input_1(wire_97), .Input_2(wire_29), .Output(wire_1));
  mand # (.UUID(64'd1055636189021926738 ^ UUID)) mand_124 (.clk(clk), .rst(rst), .Input_1(wire_64), .Input_2(wire_29), .Output(wire_8));
  mand # (.UUID(64'd3603338431621519469 ^ UUID)) mand_125 (.clk(clk), .rst(rst), .Input_1(wire_50), .Input_2(wire_29), .Output(wire_74));
  OnOrOff # (.UUID(64'd2326604957341175433 ^ UUID)) OnOrOff_126 (.clk(clk), .rst(rst), .Input(wire_20), .Output(wire_29_0));
  _99z_Counterz_Manual # (.UUID(64'd1622372112810930977 ^ UUID)) _99z_Counterz_Manual_127 (.clk(clk), .rst(rst), .Manual_Incrment(wire_105), .Out(wire_88), .Increment(wire_106));
  _99z_Counterz_Manual # (.UUID(64'd436698719286378264 ^ UUID)) _99z_Counterz_Manual_128 (.clk(clk), .rst(rst), .Manual_Incrment(wire_27), .Out(wire_80), .Increment(wire_105));
  flippedzm64bzmswitch # (.UUID(64'd3953824495697847095 ^ UUID)) flippedzm64bzmswitch_129 (.clk(clk), .rst(rst), .Input_1(wire_107), .Input_2(wire_13), .Output(wire_98));
  OnOrOff # (.UUID(64'd1722073530503975284 ^ UUID)) OnOrOff_130 (.clk(clk), .rst(rst), .Input(wire_62), .Output(wire_40_0));
  OnOrOff # (.UUID(64'd206339419552634729 ^ UUID)) OnOrOff_131 (.clk(clk), .rst(rst), .Input(wire_81), .Output(wire_7_0));
  OnOrOff # (.UUID(64'd1737851237083279124 ^ UUID)) OnOrOff_132 (.clk(clk), .rst(rst), .Input(wire_100), .Output(wire_7_1));
  flippedzm64bzmswitch # (.UUID(64'd356768830879435446 ^ UUID)) flippedzm64bzmswitch_133 (.clk(clk), .rst(rst), .Input_1(wire_36), .Input_2(wire_13), .Output(wire_9_0));
  rSwitch # (.UUID(64'd967608646389528694 ^ UUID)) rSwitch_134 (.clk(clk), .rst(rst), .Input(wire_84), .Enable(wire_13), .Output(wire_40_1));
  rSwitch # (.UUID(64'd4366678866059463544 ^ UUID)) rSwitch_135 (.clk(clk), .rst(rst), .Input(wire_29), .Enable(wire_13), .Output(wire_89));
  jump # (.UUID(64'd3373719407645708689 ^ UUID)) jump_136 (.clk(clk), .rst(rst), .Input(wire_2), .Output(wire_84));
  jump64b # (.UUID(64'd899973515945511666 ^ UUID)) jump64b_137 (.clk(clk), .rst(rst), .Input(wire_4), .Output(wire_107));
  jump64b # (.UUID(64'd2123588842821160881 ^ UUID)) jump64b_138 (.clk(clk), .rst(rst), .Input(wire_19), .Output(wire_36));
  _64zmany # (.UUID(64'd1931968964033189129 ^ UUID)) _64zmany_139 (.clk(clk), .rst(rst), .Input(wire_5), .Output(wire_48));
  OnOrOff # (.UUID(64'd4135007685282140821 ^ UUID)) OnOrOff_140 (.clk(clk), .rst(rst), .Input(wire_91), .Output(wire_78_0));

  wire [63:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_2_0;
  wire [0:0] wire_2_1;
  assign wire_2 = wire_2_0|wire_2_1;
  wire [0:0] wire_3;
  wire [63:0] wire_4;
  wire [63:0] wire_4_0;
  wire [63:0] wire_4_1;
  assign wire_4 = wire_4_0|wire_4_1;
  wire [63:0] wire_5;
  wire [7:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_7_0;
  wire [0:0] wire_7_1;
  assign wire_7 = wire_7_0|wire_7_1;
  wire [0:0] wire_8;
  wire [63:0] wire_9;
  wire [63:0] wire_9_0;
  wire [63:0] wire_9_1;
  assign wire_9 = wire_9_0|wire_9_1;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [63:0] wire_12;
  wire [0:0] wire_13;
  wire [63:0] wire_14;
  wire [0:0] wire_15;
  wire [63:0] wire_16;
  wire [0:0] wire_17;
  wire [63:0] wire_18;
  wire [63:0] wire_19;
  wire [63:0] wire_19_0;
  wire [63:0] wire_19_1;
  wire [63:0] wire_19_2;
  wire [63:0] wire_19_3;
  assign wire_19 = wire_19_0|wire_19_1|wire_19_2|wire_19_3;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [63:0] wire_22;
  wire [7:0] wire_23;
  wire [7:0] wire_23_0;
  wire [7:0] wire_23_1;
  wire [7:0] wire_23_2;
  assign wire_23 = wire_23_0|wire_23_1|wire_23_2;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_29_0;
  wire [0:0] wire_29_1;
  wire [0:0] wire_29_2;
  assign wire_29 = wire_29_0|wire_29_1|wire_29_2;
  wire [63:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [63:0] wire_33;
  wire [0:0] wire_34;
  wire [63:0] wire_35;
  wire [63:0] wire_35_0;
  wire [63:0] wire_35_1;
  wire [63:0] wire_35_2;
  wire [63:0] wire_35_3;
  wire [63:0] wire_35_4;
  wire [63:0] wire_35_5;
  assign wire_35 = wire_35_0|wire_35_1|wire_35_2|wire_35_3|wire_35_4|wire_35_5;
  wire [63:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_38_0;
  wire [0:0] wire_38_1;
  assign wire_38 = wire_38_0|wire_38_1;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_40_0;
  wire [0:0] wire_40_1;
  assign wire_40 = wire_40_0|wire_40_1;
  wire [63:0] wire_41;
  wire [0:0] wire_42;
  wire [63:0] wire_43;
  wire [63:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [63:0] wire_47;
  wire [63:0] wire_47_0;
  wire [63:0] wire_47_1;
  assign wire_47 = wire_47_0|wire_47_1;
  wire [0:0] wire_48;
  wire [63:0] wire_49;
  wire [0:0] wire_50;
  wire [63:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [7:0] wire_54;
  wire [0:0] wire_55;
  wire [63:0] wire_56;
  wire [63:0] wire_57;
  wire [63:0] wire_58;
  wire [63:0] wire_59;
  wire [63:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [63:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [63:0] wire_66;
  wire [63:0] wire_67;
  wire [63:0] wire_67_0;
  wire [63:0] wire_67_1;
  assign wire_67 = wire_67_0|wire_67_1;
  wire [0:0] wire_68;
  wire [63:0] wire_69;
  wire [63:0] wire_70;
  wire [63:0] wire_71;
  wire [0:0] wire_72;
  assign wire_72 = 0;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [63:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_78_0;
  wire [0:0] wire_78_1;
  assign wire_78 = wire_78_0|wire_78_1;
  wire [0:0] wire_79;
  wire [7:0] wire_80;
  wire [0:0] wire_81;
  wire [63:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [7:0] wire_88;
  wire [0:0] wire_89;
  wire [63:0] wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  wire [63:0] wire_93;
  wire [63:0] wire_94;
  wire [0:0] wire_95;
  wire [0:0] wire_96;
  wire [0:0] wire_97;
  wire [63:0] wire_98;
  wire [7:0] wire_99;
  wire [0:0] wire_100;
  wire [63:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [0:0] wire_106;
  wire [63:0] wire_107;
  wire [0:0] wire_108;
  wire [0:0] wire_109;
  wire [7:0] wire_110;

endmodule
