module _64zmany (clk, rst, Input, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [63:0] Input;
  output  wire [0:0] Output;

  TC_Splitter64 # (.UUID(64'd4125071985560356186 ^ UUID)) Splitter64_0 (.in(wire_9), .out0(wire_2), .out1(wire_1), .out2(wire_7), .out3(wire_3), .out4(wire_5), .out5(wire_6), .out6(wire_4), .out7(wire_8));
  _8zmany # (.UUID(64'd3464223514687233175 ^ UUID)) _8zmany_1 (.clk(clk), .rst(rst), .Input(wire_2), .Output(wire_0_5));
  _8zmany # (.UUID(64'd4137999141185627173 ^ UUID)) _8zmany_2 (.clk(clk), .rst(rst), .Input(wire_1), .Output(wire_0_3));
  _8zmany # (.UUID(64'd3788585425594785226 ^ UUID)) _8zmany_3 (.clk(clk), .rst(rst), .Input(wire_7), .Output(wire_0_0));
  _8zmany # (.UUID(64'd4259720684948900868 ^ UUID)) _8zmany_4 (.clk(clk), .rst(rst), .Input(wire_3), .Output(wire_0_1));
  _8zmany # (.UUID(64'd2794389762005023904 ^ UUID)) _8zmany_5 (.clk(clk), .rst(rst), .Input(wire_5), .Output(wire_0_2));
  _8zmany # (.UUID(64'd3111178828825728487 ^ UUID)) _8zmany_6 (.clk(clk), .rst(rst), .Input(wire_6), .Output(wire_0_4));
  _8zmany # (.UUID(64'd4522525665121392228 ^ UUID)) _8zmany_7 (.clk(clk), .rst(rst), .Input(wire_4), .Output(wire_0_6));
  _8zmany # (.UUID(64'd3883398377266044185 ^ UUID)) _8zmany_8 (.clk(clk), .rst(rst), .Input(wire_8), .Output(wire_0_7));
  TC_Switch # (.UUID(64'd666363699208919671 ^ UUID), .BIT_WIDTH(64'd1)) Output1z_9 (.en(wire_0), .in(wire_0), .out(Output));

  wire [0:0] wire_0;
  wire [0:0] wire_0_0;
  wire [0:0] wire_0_1;
  wire [0:0] wire_0_2;
  wire [0:0] wire_0_3;
  wire [0:0] wire_0_4;
  wire [0:0] wire_0_5;
  wire [0:0] wire_0_6;
  wire [0:0] wire_0_7;
  assign wire_0 = wire_0_0|wire_0_1|wire_0_2|wire_0_3|wire_0_4|wire_0_5|wire_0_6|wire_0_7;
  wire [7:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_3;
  wire [7:0] wire_4;
  wire [7:0] wire_5;
  wire [7:0] wire_6;
  wire [7:0] wire_7;
  wire [7:0] wire_8;
  wire [63:0] wire_9;
  assign wire_9 = Input;

endmodule
