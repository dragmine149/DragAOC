module _99z_Counterz_Manual (clk, rst, Manual_Incrment, Out, Increment);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] Manual_Incrment;
  output  wire [7:0] Out;
  output  wire [0:0] Increment;

  TC_DelayLine # (.UUID(64'd34289904509194689 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_0 (.clk(clk), .rst(rst), .in(wire_3), .out(wire_36));
  TC_DelayLine # (.UUID(64'd4069358971013078268 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_1 (.clk(clk), .rst(rst), .in(wire_2), .out(wire_39));
  TC_DelayLine # (.UUID(64'd738497110400040061 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_2 (.clk(clk), .rst(rst), .in(wire_9), .out(wire_34));
  TC_DelayLine # (.UUID(64'd4346959709694729258 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_3 (.clk(clk), .rst(rst), .in(wire_17), .out(wire_22));
  TC_DelayLine # (.UUID(64'd1725319397674810636 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_4 (.clk(clk), .rst(rst), .in(wire_21), .out(wire_43));
  TC_DelayLine # (.UUID(64'd47721268601486515 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_5 (.clk(clk), .rst(rst), .in(wire_1), .out(wire_32));
  TC_DelayLine # (.UUID(64'd3592910104999865036 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_6 (.clk(clk), .rst(rst), .in(wire_13), .out(wire_29));
  TC_And3 # (.UUID(64'd65592815809949785 ^ UUID), .BIT_WIDTH(64'd1)) And3_7 (.in0(wire_4), .in1(wire_10), .in2(wire_16), .out(wire_19));
  TC_And # (.UUID(64'd3024611099915004594 ^ UUID), .BIT_WIDTH(64'd1)) And_8 (.in0(wire_19), .in1(wire_5), .out(wire_6));
  TC_Not # (.UUID(64'd3161378712174442265 ^ UUID), .BIT_WIDTH(64'd1)) Not_9 (.in(wire_5), .out(wire_44));
  TC_Not # (.UUID(64'd2327727388980912896 ^ UUID), .BIT_WIDTH(64'd1)) Not_10 (.in(wire_45), .out(wire_0));
  _7bitz_Maker # (.UUID(64'd1696673967891224118 ^ UUID)) _7bitz_Maker_11 (.clk(clk), .rst(rst), .\1 (wire_43), .\2 (wire_22), .\4 (wire_34), .\8 (wire_39), .\16 (wire_36), .\32 (wire_29), .\64 (wire_32), .Output(wire_24));
  _7bitz_Seperator # (.UUID(64'd4251408542555170009 ^ UUID)) _7bitz_Seperator_12 (.clk(clk), .rst(rst), .Input(wire_24), .\1 (wire_5), .\2 (wire_16), .\4 (wire_23), .\8 (wire_18), .\16 (wire_14), .\32 (wire_10), .\64 (wire_4));
  xorandoutputswitchz_NC # (.UUID(64'd4298636058826096025 ^ UUID)) xorandoutputswitchz_NC_13 (.clk(clk), .rst(rst), .Bit(wire_4), .Carry(wire_35), .Overrite_bit(1'd0), .Overite(wire_42), .Output(wire_30));
  xorandoutputswitch # (.UUID(64'd1586845958422630920 ^ UUID)) xorandoutputswitch_14 (.clk(clk), .rst(rst), .Bit(wire_10), .Carry(wire_26), .Overrite_bit(1'd0), .Overite(wire_11), .Overrite(wire_42), .And(wire_35), .Output(wire_41));
  xorandoutputswitch # (.UUID(64'd1521851550400027753 ^ UUID)) xorandoutputswitch_15 (.clk(clk), .rst(rst), .Bit(wire_14), .Carry(wire_37), .Overrite_bit(1'd0), .Overite(wire_12), .Overrite(wire_11), .And(wire_26), .Output(wire_46));
  xorandoutputswitch # (.UUID(64'd1489539927334991040 ^ UUID)) xorandoutputswitch_16 (.clk(clk), .rst(rst), .Bit(wire_18), .Carry(wire_28), .Overrite_bit(1'd0), .Overite(wire_33), .Overrite(wire_12), .And(wire_37), .Output(wire_7));
  xorandoutputswitch # (.UUID(64'd583007522798265788 ^ UUID)) xorandoutputswitch_17 (.clk(clk), .rst(rst), .Bit(wire_23), .Carry(wire_38), .Overrite_bit(1'd0), .Overite(wire_25), .Overrite(wire_33), .And(wire_28), .Output(wire_31));
  xorandoutputswitch # (.UUID(64'd1496681166144823165 ^ UUID)) xorandoutputswitch_18 (.clk(clk), .rst(rst), .Bit(wire_16), .Carry(wire_5), .Overrite_bit(1'd0), .Overite(wire_6), .Overrite(wire_25), .And(wire_38), .Output(wire_20));
  outputswitch # (.UUID(64'd1939714350299288130 ^ UUID)) outputswitch_19 (.clk(clk), .rst(rst), .Input_A(wire_4), .Input_B(wire_30), .Path(wire_0), .Output(wire_1));
  outputswitch # (.UUID(64'd1200188231228578026 ^ UUID)) outputswitch_20 (.clk(clk), .rst(rst), .Input_A(wire_10), .Input_B(wire_41), .Path(wire_0), .Output(wire_13));
  outputswitch # (.UUID(64'd2099594080562067651 ^ UUID)) outputswitch_21 (.clk(clk), .rst(rst), .Input_A(wire_14), .Input_B(wire_46), .Path(wire_0), .Output(wire_3));
  outputswitch # (.UUID(64'd813194914662741333 ^ UUID)) outputswitch_22 (.clk(clk), .rst(rst), .Input_A(wire_18), .Input_B(wire_7), .Path(wire_0), .Output(wire_2));
  outputswitch # (.UUID(64'd823390921480707477 ^ UUID)) outputswitch_23 (.clk(clk), .rst(rst), .Input_A(wire_23), .Input_B(wire_31), .Path(wire_0), .Output(wire_9));
  outputswitch # (.UUID(64'd2128035273330340028 ^ UUID)) outputswitch_24 (.clk(clk), .rst(rst), .Input_A(wire_16), .Input_B(wire_20), .Path(wire_0), .Output(wire_17));
  outputswitch # (.UUID(64'd4438166323728123426 ^ UUID)) outputswitch_25 (.clk(clk), .rst(rst), .Input_A(wire_5), .Input_B(wire_44), .Path(wire_0), .Output(wire_21));
  _7bitz_Maker # (.UUID(64'd1681064825966949001 ^ UUID)) _7bitz_Maker_26 (.clk(clk), .rst(rst), .\1 (wire_1), .\2 (wire_13), .\4 (wire_3), .\8 (wire_2), .\16 (wire_9), .\32 (wire_17), .\64 (wire_21), .Output(wire_40));
  _8zmany # (.UUID(64'd3755729894865580756 ^ UUID)) _8zmany_27 (.clk(clk), .rst(rst), .Input(wire_40), .Output(wire_8));
  mand # (.UUID(64'd2808018554483345532 ^ UUID)) mand_28 (.clk(clk), .rst(rst), .Input_1(wire_15), .Input_2(wire_6), .Output(wire_27));
  TC_Not # (.UUID(64'd190037023794496435 ^ UUID), .BIT_WIDTH(64'd1)) Not_29 (.in(wire_8), .out(wire_15));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [0:0] wire_11;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [7:0] wire_24;
  assign Out = wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  assign Increment = wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [7:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  assign wire_45 = Manual_Incrment;
  wire [0:0] wire_46;

endmodule
