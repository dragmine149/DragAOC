module Day3Part1z_Attempt3 (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_FileLoader # (.UUID(64'd670867910265240022 ^ UUID), .DEFAULT_FILE_NAME("day3")) FileLoader_0 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_0), .out(wire_8_0));
  TC_Constant # (.UUID(64'd3936697611034503221 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_1 (.out());
  TC_FileLoader # (.UUID(64'd1471818332144234541 ^ UUID), .DEFAULT_FILE_NAME("day3_test_1")) FileLoader_2 (.clk(clk), .rst(rst), .en(wire_59), .address(wire_0), .out(wire_8_1));
  TC_Constant # (.UUID(64'd3499631194368056916 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_3 (.out(wire_59));
  TC_Constant # (.UUID(64'd2232736622141656856 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_4 (.out());
  TC_Constant # (.UUID(64'd1981730186504267880 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_5 (.out());
  TC_Constant # (.UUID(64'd1021525384996764303 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_6 (.out());
  TC_Constant # (.UUID(64'd2233006607170672073 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_7 (.out());
  TC_Constant # (.UUID(64'd2545521340778047509 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_8 (.out());
  TC_Constant # (.UUID(64'd106938163112223798 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_9 (.out());
  TC_Constant # (.UUID(64'd4318802647083067959 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_10 (.out());
  TC_Constant # (.UUID(64'd1130820721428926793 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_11 (.out());
  TC_Constant # (.UUID(64'd291644535782022576 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_12 (.out());
  TC_Constant # (.UUID(64'd4226570772319391860 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_13 (.out());
  TC_Constant # (.UUID(64'd2621130069460615979 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_14 (.out());
  TC_Constant # (.UUID(64'd810286633950345646 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_15 (.out());
  TC_Constant # (.UUID(64'd154484762821244521 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_16 (.out());
  TC_Constant # (.UUID(64'd1293101044721837465 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_17 (.out());
  TC_Constant # (.UUID(64'd1919304839526120989 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFFFFFFFFFFFFFFFF)) Constant64_18 (.out(wire_42));
  TC_Add # (.UUID(64'd539826787227496491 ^ UUID), .BIT_WIDTH(64'd64)) Add64_19 (.in0(wire_73), .in1(wire_23), .ci(1'd0), .out(wire_26), .co());
  TC_DelayLine # (.UUID(64'd1121378025258459254 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_20 (.clk(clk), .rst(rst), .in(wire_26), .out(wire_23));
  TC_Mux # (.UUID(64'd400526689135511509 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_21 (.sel(wire_39), .in0(wire_42), .in1(wire_23), .out(wire_0));
  TC_Switch # (.UUID(64'd3750085722990771933 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_22 (.en(wire_39), .in({{56{1'b0}}, wire_21 }), .out(wire_73));
  TC_Equal # (.UUID(64'd1006503156420949217 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_23 (.in0(wire_23), .in1(wire_7), .out(wire_32));
  TC_And3 # (.UUID(64'd330147788875224171 ^ UUID), .BIT_WIDTH(64'd1)) And3_24 (.in0(wire_54), .in1(wire_56), .in2(wire_77), .out(wire_39));
  TC_Not # (.UUID(64'd285764211932754545 ^ UUID), .BIT_WIDTH(64'd1)) Not_25 (.in(wire_32), .out(wire_77));
  TC_Counter # (.UUID(64'd1078548748747073918 ^ UUID), .BIT_WIDTH(64'd32), .count(32'd1)) Counter32_26 (.clk(clk), .rst(rst), .save(wire_27), .in(wire_65), .out(wire_22));
  TC_Ram # (.UUID(64'd889594913348838705 ^ UUID), .WORD_WIDTH(64'd32), .WORD_COUNT(64'd384)) Ram_27 (.clk(clk), .rst(rst), .load(wire_50[0:0]), .save(wire_47), .address(wire_22), .in0({{32{1'b0}}, wire_3 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_33), .out1(), .out2(), .out3());
  TC_Splitter32 # (.UUID(64'd4035469326953262772 ^ UUID)) Splitter32_28 (.in(wire_81), .out0(wire_14), .out1(wire_60), .out2(wire_57), .out3(wire_9));
  TC_Maker16 # (.UUID(64'd3928271251860206036 ^ UUID)) Maker16_29 (.in0(wire_14), .in1(wire_60), .out(wire_20));
  TC_Maker16 # (.UUID(64'd3642668000385795629 ^ UUID)) Maker16_30 (.in0(wire_57), .in1(wire_9), .out(wire_83));
  TC_DelayLine # (.UUID(64'd1069740274028324431 ^ UUID), .BIT_WIDTH(64'd32)) DelayLine32_31 (.clk(clk), .rst(rst), .in(wire_71), .out(wire_19));
  TC_Mux # (.UUID(64'd1933241523835954014 ^ UUID), .BIT_WIDTH(64'd32)) Mux32_32 (.sel(wire_35), .in0(wire_19), .in1({{24{1'b0}}, wire_43 }), .out(wire_66));
  TC_Mux # (.UUID(64'd3591417222352229250 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_33 (.sel(wire_6), .in0(wire_19[7:0]), .in1(wire_28[7:0]), .out(wire_43));
  TC_LessI # (.UUID(64'd4164544218120390221 ^ UUID), .BIT_WIDTH(64'd32)) LessI32_34 (.in0(wire_28), .in1(wire_19), .out(wire_6));
  TC_Constant # (.UUID(64'd896447414079347299 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h7FFFFFFF)) Constant32_35 (.out(wire_78));
  TC_Constant # (.UUID(64'd503246965407474427 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_36 (.out(wire_29));
  TC_DelayLine # (.UUID(64'd3658476492014616617 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_37 (.clk(clk), .rst(rst), .in(wire_29), .out(wire_2));
  TC_Switch # (.UUID(64'd3341655025280185596 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_38 (.en(wire_2), .in(wire_66), .out(wire_71_1));
  TC_Switch # (.UUID(64'd3193310534451515930 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_39 (.en(wire_31), .in(wire_78), .out(wire_71_0));
  TC_Switch # (.UUID(64'd317804265825901077 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_40 (.en(wire_68), .in(wire_29), .out(wire_31));
  TC_Not # (.UUID(64'd919022448505067535 ^ UUID), .BIT_WIDTH(64'd1)) Not_41 (.in(wire_2), .out(wire_68));
  TC_DelayLine # (.UUID(64'd600003832322404005 ^ UUID), .BIT_WIDTH(64'd32)) DelayLine32_42 (.clk(clk), .rst(rst), .in(wire_33[31:0]), .out(wire_30));
  TC_Splitter32 # (.UUID(64'd4155479272641838016 ^ UUID)) Splitter32_43 (.in(wire_79), .out0(wire_18), .out1(wire_1), .out2(wire_64), .out3(wire_69));
  TC_Maker16 # (.UUID(64'd1243116669575388859 ^ UUID)) Maker16_44 (.in0(wire_18), .in1(wire_1), .out(wire_44));
  TC_Maker16 # (.UUID(64'd1497221609392710490 ^ UUID)) Maker16_45 (.in0(wire_64), .in1(wire_69), .out(wire_63));
  TC_Splitter32 # (.UUID(64'd1230841868525626631 ^ UUID)) Splitter32_46 (.in(wire_5), .out0(wire_17), .out1(wire_38), .out2(wire_67), .out3(wire_75));
  TC_Maker16 # (.UUID(64'd1644724077454726226 ^ UUID)) Maker16_47 (.in0(wire_17), .in1(wire_38), .out(wire_37));
  TC_Maker16 # (.UUID(64'd2152189888456059487 ^ UUID)) Maker16_48 (.in0(wire_67), .in1(wire_75), .out(wire_41));
  TC_Splitter32 # (.UUID(64'd4418466857278764279 ^ UUID)) Splitter32_49 (.in(wire_33[31:0]), .out0(wire_52), .out1(wire_10), .out2(wire_45), .out3(wire_62));
  TC_Maker16 # (.UUID(64'd3349853774350948360 ^ UUID)) Maker16_50 (.in0(wire_52), .in1(wire_10), .out(wire_82));
  TC_Maker16 # (.UUID(64'd2883050298416608739 ^ UUID)) Maker16_51 (.in0(wire_45), .in1(wire_62), .out(wire_46));
  TC_Splitter32 # (.UUID(64'd230254807600720706 ^ UUID)) Splitter32_52 (.in(wire_30), .out0(wire_36), .out1(wire_48), .out2(wire_72), .out3(wire_16));
  TC_Maker16 # (.UUID(64'd2484952494794539159 ^ UUID)) Maker16_53 (.in0(wire_36), .in1(wire_48), .out(wire_25));
  TC_Maker16 # (.UUID(64'd1925151316157446563 ^ UUID)) Maker16_54 (.in0(wire_72), .in1(wire_16), .out(wire_15));
  TC_Not # (.UUID(64'd3539672329771887091 ^ UUID), .BIT_WIDTH(64'd1)) Not_55 (.in(wire_34), .out(wire_40));
  TC_Mux # (.UUID(64'd869346753072203086 ^ UUID), .BIT_WIDTH(64'd32)) Mux32_56 (.sel(wire_27), .in0(wire_22), .in1(32'd0), .out(wire_65));
  TC_Not # (.UUID(64'd1498694609800071896 ^ UUID), .BIT_WIDTH(64'd1)) Not_57 (.in(wire_76), .out(wire_11));
  TC_Not # (.UUID(64'd1524827408234024151 ^ UUID), .BIT_WIDTH(64'd1)) Not_58 (.in(wire_49), .out(wire_47));
  TC_And3 # (.UUID(64'd3042879754477079505 ^ UUID), .BIT_WIDTH(64'd1)) And3_59 (.in0(wire_40), .in1(wire_51), .in2(wire_53), .out(wire_76));
  TC_Equal # (.UUID(64'd3161989386235867289 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_60 (.in0(wire_22), .in1(wire_55[31:0]), .out(wire_24));
  TC_Switch # (.UUID(64'd948381973252070923 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_61 (.en(wire_34), .in(wire_22), .out(wire_70));
  TC_Not # (.UUID(64'd1674548457943997484 ^ UUID), .BIT_WIDTH(64'd1)) Not_62 (.in(wire_13), .out(wire_53));
  TC_And # (.UUID(64'd2893488111660484409 ^ UUID), .BIT_WIDTH(64'd1)) And_63 (.in0(wire_24), .in1(wire_4), .out(wire_13));
  TC_Halt # (.UUID(64'd1474802306642119463 ^ UUID), .HALT_MESSAGE("End of file reached!")) Halt_64 (.clk(clk), .rst(rst), .en(wire_74));
  TC_DelayLine # (.UUID(64'd476274355105221649 ^ UUID), .BIT_WIDTH(64'd32)) DelayLine32_65 (.clk(clk), .rst(rst), .in(wire_3), .out(wire_80));
  TC_Halt # (.UUID(64'd3727559317572521050 ^ UUID), .HALT_MESSAGE("Found crossing")) Halt_66 (.clk(clk), .rst(rst), .en(1'd0));
  TC_And3 # (.UUID(64'd3134744527415087055 ^ UUID), .BIT_WIDTH(64'd1)) And3_67 (.in0(wire_56), .in1(wire_13), .in2(wire_32), .out(wire_74));
  TC_FileLoader # (.UUID(64'd3429124062269983960 ^ UUID), .DEFAULT_FILE_NAME("day3_test_2")) FileLoader_68 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_0), .out(wire_8_2));
  TC_FileLoader # (.UUID(64'd1473616339079632962 ^ UUID), .DEFAULT_FILE_NAME("day3_test_3")) FileLoader_69 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_0), .out(wire_8_3));
  InputMananger # (.UUID(64'd280349663464583758 ^ UUID)) InputMananger_70 (.clk(clk), .rst(rst), .Main_8b(wire_8), .Offset(wire_21), .Output(wire_12), .NewLine(wire_34));
  QuickSave # (.UUID(64'd3964331221245691836 ^ UUID)) QuickSave_71 (.clk(clk), .rst(rst), .Value(wire_8), .\Number_(stored) (wire_7), .\Saved?_1 (wire_56), .\Saved?_2 (wire_51));
  ManhattanDistance # (.UUID(64'd4534475870914388036 ^ UUID)) ManhattanDistance_72 (.clk(clk), .rst(rst), .Y(wire_83), .X(wire_20), .Output(wire_28));
  CellRotator # (.UUID(64'd2988738449177159528 ^ UUID)) CellRotator_73 (.clk(clk), .rst(rst), .Input(wire_58), .Tick(wire_13), .Pos_2(wire_5), .Pos_1(wire_79), .Written());
  QuickSave # (.UUID(64'd3551179199781681902 ^ UUID)) QuickSave_74 (.clk(clk), .rst(rst), .Value({{63{1'b0}}, wire_34 }), .\Number_(stored) (wire_50), .\Saved?_1 (wire_49), .\Saved?_2 ());
  OnOrOff # (.UUID(64'd2880407376120648954 ^ UUID)) OnOrOff_75 (.clk(clk), .rst(rst), .Input(wire_11), .Output(wire_27));
  QuickSave # (.UUID(64'd4013860832325939171 ^ UUID)) QuickSave_76 (.clk(clk), .rst(rst), .Value({{32{1'b0}}, wire_70 }), .\Number_(stored) (wire_55), .\Saved?_1 (wire_4), .\Saved?_2 ());
  OnOrOff # (.UUID(64'd685402883028759750 ^ UUID)) OnOrOff_77 (.clk(clk), .rst(rst), .Input(wire_47), .Output(wire_54_0));
  OnOrOff # (.UUID(64'd2586521289870388092 ^ UUID)) OnOrOff_78 (.clk(clk), .rst(rst), .Input(wire_13), .Output(wire_54_1));
  PositionAdder # (.UUID(64'd4180759426517963882 ^ UUID)) PositionAdder_79 (.clk(clk), .rst(rst), .Current_Position(wire_80), .Move(wire_12), .overflow(wire_61), .New_Position(wire_3));
  PositionAdder # (.UUID(64'd3058909452894868054 ^ UUID)) PositionAdder_80 (.clk(clk), .rst(rst), .Current_Position(wire_5), .Move(wire_12), .overflow(), .New_Position(wire_58));
  LineCrosserz_3 # (.UUID(64'd3547560156308371360 ^ UUID)) LineCrosserz_3_81 (.clk(clk), .rst(rst), .Input_1(wire_5), .Input_2(wire_79), .Input_3(wire_33[31:0]), .Input_4(wire_30), .Output_1(wire_35), .Output_2(wire_81));
  TC_Halt # (.UUID(64'd2886596719389344914 ^ UUID), .HALT_MESSAGE("Adder overflow! (PositionAdder)")) Halt_82 (.clk(clk), .rst(rst), .en(wire_61));

  wire [63:0] wire_0;
  wire [7:0] wire_1;
  wire [0:0] wire_2;
  wire [31:0] wire_3;
  wire [0:0] wire_4;
  wire [31:0] wire_5;
  wire [0:0] wire_6;
  wire [63:0] wire_7;
  wire [63:0] wire_8;
  wire [63:0] wire_8_0;
  wire [63:0] wire_8_1;
  wire [63:0] wire_8_2;
  wire [63:0] wire_8_3;
  assign wire_8 = wire_8_0|wire_8_1|wire_8_2|wire_8_3;
  wire [7:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [31:0] wire_12;
  wire [0:0] wire_13;
  wire [7:0] wire_14;
  wire [15:0] wire_15;
  wire [7:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_18;
  wire [31:0] wire_19;
  wire [15:0] wire_20;
  wire [7:0] wire_21;
  wire [31:0] wire_22;
  wire [63:0] wire_23;
  wire [0:0] wire_24;
  wire [15:0] wire_25;
  wire [63:0] wire_26;
  wire [0:0] wire_27;
  wire [31:0] wire_28;
  wire [0:0] wire_29;
  wire [31:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [63:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [7:0] wire_36;
  wire [15:0] wire_37;
  wire [7:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [15:0] wire_41;
  wire [63:0] wire_42;
  wire [7:0] wire_43;
  wire [15:0] wire_44;
  wire [7:0] wire_45;
  wire [15:0] wire_46;
  wire [0:0] wire_47;
  wire [7:0] wire_48;
  wire [0:0] wire_49;
  wire [63:0] wire_50;
  wire [0:0] wire_51;
  wire [7:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_54_0;
  wire [0:0] wire_54_1;
  assign wire_54 = wire_54_0|wire_54_1;
  wire [63:0] wire_55;
  wire [0:0] wire_56;
  wire [7:0] wire_57;
  wire [31:0] wire_58;
  wire [0:0] wire_59;
  wire [7:0] wire_60;
  wire [0:0] wire_61;
  wire [7:0] wire_62;
  wire [15:0] wire_63;
  wire [7:0] wire_64;
  wire [31:0] wire_65;
  wire [31:0] wire_66;
  wire [7:0] wire_67;
  wire [0:0] wire_68;
  wire [7:0] wire_69;
  wire [31:0] wire_70;
  wire [31:0] wire_71;
  wire [31:0] wire_71_0;
  wire [31:0] wire_71_1;
  assign wire_71 = wire_71_0|wire_71_1;
  wire [7:0] wire_72;
  wire [63:0] wire_73;
  wire [0:0] wire_74;
  wire [7:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [31:0] wire_78;
  wire [31:0] wire_79;
  wire [31:0] wire_80;
  wire [31:0] wire_81;
  wire [15:0] wire_82;
  wire [15:0] wire_83;

endmodule
