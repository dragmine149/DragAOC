module LineCrosserz_3 (clk, rst, L2End, L2Start, L1End, L1Start, Intercection, Point_of_Interce, \StepCount_(r) );
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [63:0] L2End;
  input  wire [63:0] L2Start;
  input  wire [63:0] L1End;
  input  wire [63:0] L1Start;
  output  wire [0:0] Intercection;
  output  wire [63:0] Point_of_Interce;
  output  wire [31:0] \StepCount_(r) ;

  TC_Switch # (.UUID(64'd29451040430517838 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_0 (.en(wire_7), .in(wire_39), .out(wire_13));
  TC_Not # (.UUID(64'd380166382871947097 ^ UUID), .BIT_WIDTH(64'd1)) Not_1 (.in(wire_27), .out(wire_7));
  TC_Switch # (.UUID(64'd3821448631046911694 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_2 (.en(wire_38), .in(wire_27), .out(wire_1));
  TC_Not # (.UUID(64'd569669821514979918 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_13), .out(wire_38));
  TC_And3 # (.UUID(64'd1658388512215494880 ^ UUID), .BIT_WIDTH(64'd1)) And3_4 (.in0(wire_31), .in1(wire_42), .in2(wire_29), .out(wire_15));
  TC_Equal # (.UUID(64'd1462953451613577458 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_5 (.in0(wire_0), .in1(wire_18), .out(wire_4));
  TC_Equal # (.UUID(64'd2477445908053147713 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_6 (.in0(wire_33), .in1(wire_36), .out(wire_20));
  TC_Equal # (.UUID(64'd3736993343762613191 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_7 (.in0(wire_28), .in1(wire_6), .out(wire_24));
  TC_Equal # (.UUID(64'd2800749848815207265 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_8 (.in0(wire_16), .in1(wire_14), .out(wire_40));
  TC_Switch # (.UUID(64'd1144186547777792254 ^ UUID), .BIT_WIDTH(64'd64)) Output64z_9 (.en(wire_15), .in(wire_5), .out(Point_of_Interce));
  TC_Constant # (.UUID(64'd3393676726258455498 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_10 (.out(wire_26));
  TC_Switch # (.UUID(64'd1431681702512503803 ^ UUID), .BIT_WIDTH(64'd32)) Output32z_11 (.en(wire_15), .in(wire_30), .out(\StepCount_(r) ));
  TC_Add # (.UUID(64'd2159422674975698004 ^ UUID), .BIT_WIDTH(64'd32)) Add32_12 (.in0(wire_32), .in1(wire_11), .ci(1'd0), .out(wire_30), .co());
  mand # (.UUID(64'd1966732459903081054 ^ UUID)) mand_13 (.clk(clk), .rst(rst), .Input_1(wire_4), .Input_2(wire_40), .Output(wire_27));
  mand # (.UUID(64'd1967875822324122093 ^ UUID)) mand_14 (.clk(clk), .rst(rst), .Input_1(wire_20), .Input_2(wire_24), .Output(wire_39));
  mOR # (.UUID(64'd3811154444398219071 ^ UUID)) mOR_15 (.clk(clk), .rst(rst), .Input_1(wire_13), .Input_2(wire_1), .Output(wire_42));
  mand # (.UUID(64'd2282199498514448531 ^ UUID)) mand_16 (.clk(clk), .rst(rst), .Input_1(wire_34), .Input_2(wire_37), .Output(wire_41));
  mand # (.UUID(64'd4236102916636182286 ^ UUID)) mand_17 (.clk(clk), .rst(rst), .Input_1(wire_17), .Input_2(wire_35), .Output(wire_10));
  mNOR # (.UUID(64'd1044973136834131328 ^ UUID)) mNOR_18 (.clk(clk), .rst(rst), .Input_1(wire_10), .Input_2(wire_41), .Output(wire_31));
  _64bz_toz_32b # (.UUID(64'd1160700702824551150 ^ UUID)) _64bz_toz_32b_19 (.clk(clk), .rst(rst), .Input(wire_19), .Output_1(wire_14), .Output_2(wire_6));
  _64bz_toz_32b # (.UUID(64'd4249573345702729115 ^ UUID)) _64bz_toz_32b_20 (.clk(clk), .rst(rst), .Input(wire_2), .Output_1(wire_16), .Output_2(wire_28));
  _64bz_toz_32b # (.UUID(64'd3482476773988014960 ^ UUID)) _64bz_toz_32b_21 (.clk(clk), .rst(rst), .Input(wire_25), .Output_1(wire_36), .Output_2(wire_18));
  _64bz_toz_32b # (.UUID(64'd1881820232260440322 ^ UUID)) _64bz_toz_32b_22 (.clk(clk), .rst(rst), .Input(wire_8), .Output_1(wire_33), .Output_2(wire_0));
  is0z_64b # (.UUID(64'd3522606142968185792 ^ UUID)) is0z_64b_23 (.clk(clk), .rst(rst), .Input(wire_8), .Output(wire_34));
  is0z_64b # (.UUID(64'd2383929583881890307 ^ UUID)) is0z_64b_24 (.clk(clk), .rst(rst), .Input(wire_25), .Output(wire_37));
  is0z_64b # (.UUID(64'd3448954266748536719 ^ UUID)) is0z_64b_25 (.clk(clk), .rst(rst), .Input(wire_2), .Output(wire_17));
  is0z_64b # (.UUID(64'd908196902127981698 ^ UUID)) is0z_64b_26 (.clk(clk), .rst(rst), .Input(wire_19), .Output(wire_35));
  PositionChcker # (.UUID(64'd470197739512970021 ^ UUID)) PositionChcker_27 (.clk(clk), .rst(rst), .HorizontalEnd(wire_3), .VerticalEnd(wire_9), .VerticalStart(wire_22), .HorizontalStart(wire_21), .Output_1(wire_29), .Output_2(wire_5));
  BusSwitcher # (.UUID(64'd4508613529556397755 ^ UUID)) BusSwitcher_28 (.clk(clk), .rst(rst), .Line_End(wire_25), .Line_Start(wire_8), .Option_1(wire_1), .Option_2(wire_13), .Horizontal_End(wire_3_1), .Horizontal_Start(wire_21_0), .Vertical_End(wire_9_1), .Vertical_Start(wire_22_1));
  BusSwitcher # (.UUID(64'd1656550384719575395 ^ UUID)) BusSwitcher_29 (.clk(clk), .rst(rst), .Line_End(wire_19), .Line_Start(wire_2), .Option_1(wire_13), .Option_2(wire_1), .Horizontal_End(wire_3_0), .Horizontal_Start(wire_21_1), .Vertical_End(wire_9_0), .Vertical_Start(wire_22_0));
  ReverseSteps # (.UUID(64'd3016120253923149437 ^ UUID)) ReverseSteps_30 (.clk(clk), .rst(rst), .LineEnd(wire_3), .InterceptPoint(wire_5), .Direction(1'd0), .StepCount(wire_12));
  ReverseSteps # (.UUID(64'd4203095323940347482 ^ UUID)) ReverseSteps_31 (.clk(clk), .rst(rst), .LineEnd(wire_9), .InterceptPoint(wire_5), .Direction(wire_26), .StepCount(wire_23));
  _32bz_ABS # (.UUID(64'd592674821184198943 ^ UUID)) _32bz_ABS_32 (.clk(clk), .rst(rst), .Input(wire_12[31:0]), .Output(wire_32));
  _32bz_ABS # (.UUID(64'd721526827469304202 ^ UUID)) _32bz_ABS_33 (.clk(clk), .rst(rst), .Input(wire_23[31:0]), .Output(wire_11));

  wire [31:0] wire_0;
  wire [0:0] wire_1;
  wire [63:0] wire_2;
  assign wire_2 = L2Start;
  wire [63:0] wire_3;
  wire [63:0] wire_3_0;
  wire [63:0] wire_3_1;
  assign wire_3 = wire_3_0|wire_3_1;
  wire [0:0] wire_4;
  wire [63:0] wire_5;
  wire [31:0] wire_6;
  wire [0:0] wire_7;
  wire [63:0] wire_8;
  assign wire_8 = L1Start;
  wire [63:0] wire_9;
  wire [63:0] wire_9_0;
  wire [63:0] wire_9_1;
  assign wire_9 = wire_9_0|wire_9_1;
  wire [0:0] wire_10;
  wire [31:0] wire_11;
  wire [63:0] wire_12;
  wire [0:0] wire_13;
  wire [31:0] wire_14;
  wire [0:0] wire_15;
  assign Intercection = wire_15;
  wire [31:0] wire_16;
  wire [0:0] wire_17;
  wire [31:0] wire_18;
  wire [63:0] wire_19;
  assign wire_19 = L2End;
  wire [0:0] wire_20;
  wire [63:0] wire_21;
  wire [63:0] wire_21_0;
  wire [63:0] wire_21_1;
  assign wire_21 = wire_21_0|wire_21_1;
  wire [63:0] wire_22;
  wire [63:0] wire_22_0;
  wire [63:0] wire_22_1;
  assign wire_22 = wire_22_0|wire_22_1;
  wire [63:0] wire_23;
  wire [0:0] wire_24;
  wire [63:0] wire_25;
  assign wire_25 = L1End;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [31:0] wire_28;
  wire [0:0] wire_29;
  wire [31:0] wire_30;
  wire [0:0] wire_31;
  wire [31:0] wire_32;
  wire [31:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [31:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;

endmodule
