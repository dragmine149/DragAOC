module PositionChcker (clk, rst, HorizontalEnd, VerticalEnd, VerticalStart, HorizontalStart, Output_1, Output_2);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [63:0] HorizontalEnd;
  input  wire [63:0] VerticalEnd;
  input  wire [63:0] VerticalStart;
  input  wire [63:0] HorizontalStart;
  output  wire [0:0] Output_1;
  output  wire [63:0] Output_2;

  TC_Maker64 # (.UUID(64'd1043128633281648890 ^ UUID)) Maker64_0 (.in0(wire_4), .in1(wire_21), .in2(wire_5), .in3(wire_1), .in4(wire_0), .in5(wire_3), .in6(wire_8), .in7(wire_22), .out(wire_23));
  TC_Splitter64 # (.UUID(64'd2780000453321243182 ^ UUID)) Splitter64_1 (.in(wire_20), .out0(wire_9), .out1(wire_45), .out2(wire_35), .out3(wire_38), .out4(), .out5(), .out6(), .out7());
  TC_Splitter64 # (.UUID(64'd4340482490135852189 ^ UUID)) Splitter64_2 (.in(wire_42), .out0(wire_10), .out1(wire_34), .out2(wire_36), .out3(wire_29), .out4(wire_0), .out5(wire_3), .out6(wire_8), .out7(wire_22));
  TC_Splitter64 # (.UUID(64'd524827928275308427 ^ UUID)) Splitter64_3 (.in(wire_26), .out0(), .out1(), .out2(), .out3(), .out4(wire_40), .out5(wire_13), .out6(wire_33), .out7(wire_24));
  TC_Splitter64 # (.UUID(64'd295433490093758283 ^ UUID)) Splitter64_4 (.in(wire_41), .out0(wire_4), .out1(wire_21), .out2(wire_5), .out3(wire_1), .out4(wire_32), .out5(wire_6), .out6(wire_27), .out7(wire_28));
  TC_Maker32 # (.UUID(64'd2951907508458143177 ^ UUID)) Maker32_5 (.in0(wire_32), .in1(wire_6), .in2(wire_27), .in3(wire_28), .out(wire_14));
  TC_Maker32 # (.UUID(64'd1903954920290057481 ^ UUID)) Maker32_6 (.in0(wire_40), .in1(wire_13), .in2(wire_33), .in3(wire_24), .out(wire_37));
  TC_Maker32 # (.UUID(64'd2975524749386368036 ^ UUID)) Maker32_7 (.in0(wire_10), .in1(wire_34), .in2(wire_36), .in3(wire_29), .out(wire_12));
  TC_Maker32 # (.UUID(64'd290392184541267702 ^ UUID)) Maker32_8 (.in0(wire_9), .in1(wire_45), .in2(wire_35), .in3(wire_38), .out(wire_47));
  TC_Maker32 # (.UUID(64'd1853444403247454946 ^ UUID)) Maker32_9 (.in0(wire_0), .in1(wire_3), .in2(wire_8), .in3(wire_22), .out(wire_19));
  TC_Maker32 # (.UUID(64'd3814693169101109449 ^ UUID)) Maker32_10 (.in0(wire_4), .in1(wire_21), .in2(wire_5), .in3(wire_1), .out(wire_2));
  TC_Switch # (.UUID(64'd4610820402517192475 ^ UUID), .BIT_WIDTH(64'd64)) Output64z_11 (.en(wire_31), .in(wire_23), .out(Output_2));
  TC_Constant # (.UUID(64'd4204772562336863462 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_12 (.out());
  mand # (.UUID(64'd4340687300676184839 ^ UUID)) mand_13 (.clk(clk), .rst(rst), .Input_1(wire_7), .Input_2(wire_18), .Output(wire_31));
  gte # (.UUID(64'd1468068711304085687 ^ UUID)) gte_14 (.clk(clk), .rst(rst), .Input_1(wire_19), .Input_2(wire_11[31:0]), .Output(wire_25));
  lte # (.UUID(64'd3067920624139790206 ^ UUID)) lte_15 (.clk(clk), .rst(rst), .Input_1(wire_19), .Input_2(wire_43[31:0]), .Output(wire_44));
  mand # (.UUID(64'd2335140900931170736 ^ UUID)) mand_16 (.clk(clk), .rst(rst), .Input_1(wire_44), .Input_2(wire_25), .Output(wire_7));
  gte # (.UUID(64'd478955746293580995 ^ UUID)) gte_17 (.clk(clk), .rst(rst), .Input_1(wire_2), .Input_2(wire_15[31:0]), .Output(wire_16));
  lte # (.UUID(64'd214932175809081470 ^ UUID)) lte_18 (.clk(clk), .rst(rst), .Input_1(wire_2), .Input_2(wire_39[31:0]), .Output(wire_46));
  mand # (.UUID(64'd300477794743194606 ^ UUID)) mand_19 (.clk(clk), .rst(rst), .Input_1(wire_46), .Input_2(wire_16), .Output(wire_18));
  minmaxz_32b # (.UUID(64'd2941986681133121684 ^ UUID)) minmaxz_32b_20 (.clk(clk), .rst(rst), .X({{32{1'b0}}, wire_14 }), .Y({{32{1'b0}}, wire_37 }), .Minimum(wire_11), .Maximum(wire_43));
  minmaxz_32b # (.UUID(64'd1487961136758229526 ^ UUID)) minmaxz_32b_21 (.clk(clk), .rst(rst), .X({{32{1'b0}}, wire_12 }), .Y({{32{1'b0}}, wire_47 }), .Minimum(wire_15), .Maximum(wire_39));
  _64bz_toz_32b # (.UUID(64'd2946613380538701206 ^ UUID)) _64bz_toz_32b_22 (.clk(clk), .rst(rst), .Input(wire_23), .Output_1(wire_17), .Output_2(wire_30));

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  wire [31:0] wire_2;
  wire [7:0] wire_3;
  wire [7:0] wire_4;
  wire [7:0] wire_5;
  wire [7:0] wire_6;
  wire [0:0] wire_7;
  wire [7:0] wire_8;
  wire [7:0] wire_9;
  wire [7:0] wire_10;
  wire [63:0] wire_11;
  wire [31:0] wire_12;
  wire [7:0] wire_13;
  wire [31:0] wire_14;
  wire [63:0] wire_15;
  wire [0:0] wire_16;
  wire [31:0] wire_17;
  wire [0:0] wire_18;
  wire [31:0] wire_19;
  wire [63:0] wire_20;
  assign wire_20 = HorizontalEnd;
  wire [7:0] wire_21;
  wire [7:0] wire_22;
  wire [63:0] wire_23;
  wire [7:0] wire_24;
  wire [0:0] wire_25;
  wire [63:0] wire_26;
  assign wire_26 = VerticalEnd;
  wire [7:0] wire_27;
  wire [7:0] wire_28;
  wire [7:0] wire_29;
  wire [31:0] wire_30;
  wire [0:0] wire_31;
  assign Output_1 = wire_31;
  wire [7:0] wire_32;
  wire [7:0] wire_33;
  wire [7:0] wire_34;
  wire [7:0] wire_35;
  wire [7:0] wire_36;
  wire [31:0] wire_37;
  wire [7:0] wire_38;
  wire [63:0] wire_39;
  wire [7:0] wire_40;
  wire [63:0] wire_41;
  assign wire_41 = VerticalStart;
  wire [63:0] wire_42;
  assign wire_42 = HorizontalStart;
  wire [63:0] wire_43;
  wire [0:0] wire_44;
  wire [7:0] wire_45;
  wire [0:0] wire_46;
  wire [31:0] wire_47;

endmodule
