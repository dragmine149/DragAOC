module Day3Part1z_Attempt3z_ZL32bZR (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_FileLoader # (.UUID(64'd670867910265240022 ^ UUID), .DEFAULT_FILE_NAME("day3")) FileLoader_0 (.clk(clk), .rst(rst), .en(wire_53), .address(wire_25), .out(wire_5_2));
  TC_Constant # (.UUID(64'd3936697611034503221 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_1 (.out(wire_53));
  TC_FileLoader # (.UUID(64'd1471818332144234541 ^ UUID), .DEFAULT_FILE_NAME("day3_test_1")) FileLoader_2 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_25), .out(wire_5_0));
  TC_Constant # (.UUID(64'd3499631194368056916 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_3 (.out());
  TC_Constant # (.UUID(64'd2232736622141656856 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_4 (.out());
  TC_Constant # (.UUID(64'd1981730186504267880 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_5 (.out());
  TC_Constant # (.UUID(64'd1021525384996764303 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_6 (.out());
  TC_Constant # (.UUID(64'd2233006607170672073 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_7 (.out());
  TC_Constant # (.UUID(64'd2545521340778047509 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_8 (.out());
  TC_Constant # (.UUID(64'd106938163112223798 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_9 (.out());
  TC_Constant # (.UUID(64'd4318802647083067959 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_10 (.out());
  TC_Constant # (.UUID(64'd1130820721428926793 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_11 (.out());
  TC_Constant # (.UUID(64'd291644535782022576 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_12 (.out());
  TC_Constant # (.UUID(64'd4226570772319391860 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_13 (.out());
  TC_Constant # (.UUID(64'd2621130069460615979 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_14 (.out());
  TC_Constant # (.UUID(64'd810286633950345646 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_15 (.out());
  TC_Constant # (.UUID(64'd154484762821244521 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_16 (.out());
  TC_Constant # (.UUID(64'd1293101044721837465 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_17 (.out());
  TC_Constant # (.UUID(64'd1919304839526120989 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFFFFFFFFFFFFFFFF)) Constant64_18 (.out(wire_35));
  TC_Add # (.UUID(64'd539826787227496491 ^ UUID), .BIT_WIDTH(64'd64)) Add64_19 (.in0(wire_45), .in1(wire_41), .ci(1'd0), .out(wire_55), .co());
  TC_DelayLine # (.UUID(64'd1121378025258459254 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_20 (.clk(clk), .rst(rst), .in(wire_55), .out(wire_41));
  TC_Mux # (.UUID(64'd400526689135511509 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_21 (.sel(wire_16), .in0(wire_35), .in1(wire_41), .out(wire_25));
  TC_Switch # (.UUID(64'd3750085722990771933 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_22 (.en(wire_16), .in({{56{1'b0}}, wire_62 }), .out(wire_45));
  TC_Equal # (.UUID(64'd1006503156420949217 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_23 (.in0(wire_41), .in1(wire_37), .out(wire_12));
  TC_And3 # (.UUID(64'd330147788875224171 ^ UUID), .BIT_WIDTH(64'd1)) And3_24 (.in0(wire_19), .in1(wire_0), .in2(wire_64), .out(wire_16));
  TC_Not # (.UUID(64'd285764211932754545 ^ UUID), .BIT_WIDTH(64'd1)) Not_25 (.in(wire_12), .out(wire_64));
  TC_Ram # (.UUID(64'd889594913348838705 ^ UUID), .WORD_WIDTH(64'd64), .WORD_COUNT(64'd512)) Ram_26 (.clk(clk), .rst(rst), .load(wire_43[0:0]), .save(wire_26), .address(wire_14), .in0(wire_18), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_22), .out1(), .out2(), .out3());
  TC_Constant # (.UUID(64'd503246965407474427 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_27 (.out(wire_60));
  TC_DelayLine # (.UUID(64'd3658476492014616617 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_28 (.clk(clk), .rst(rst), .in(wire_60), .out(wire_9));
  TC_Switch # (.UUID(64'd317804265825901077 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_29 (.en(wire_21), .in(wire_60), .out(wire_57));
  TC_Not # (.UUID(64'd919022448505067535 ^ UUID), .BIT_WIDTH(64'd1)) Not_30 (.in(wire_9), .out(wire_21));
  TC_Not # (.UUID(64'd3539672329771887091 ^ UUID), .BIT_WIDTH(64'd1)) Not_31 (.in(wire_44), .out(wire_6));
  TC_Mux # (.UUID(64'd869346753072203086 ^ UUID), .BIT_WIDTH(64'd32)) Mux32_32 (.sel(wire_24), .in0(wire_14), .in1(32'd0), .out(wire_51));
  TC_Not # (.UUID(64'd1498694609800071896 ^ UUID), .BIT_WIDTH(64'd1)) Not_33 (.in(wire_52), .out(wire_65));
  TC_Not # (.UUID(64'd1524827408234024151 ^ UUID), .BIT_WIDTH(64'd1)) Not_34 (.in(wire_47), .out(wire_26));
  TC_And3 # (.UUID(64'd3042879754477079505 ^ UUID), .BIT_WIDTH(64'd1)) And3_35 (.in0(wire_6), .in1(wire_56), .in2(wire_36), .out(wire_52));
  TC_Equal # (.UUID(64'd3161989386235867289 ^ UUID), .BIT_WIDTH(64'd32)) Equal32_36 (.in0(wire_14), .in1(wire_42[31:0]), .out(wire_48));
  TC_Switch # (.UUID(64'd948381973252070923 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_37 (.en(wire_44), .in(wire_14), .out(wire_10));
  TC_Not # (.UUID(64'd1674548457943997484 ^ UUID), .BIT_WIDTH(64'd1)) Not_38 (.in(wire_20), .out(wire_36));
  TC_And # (.UUID(64'd2893488111660484409 ^ UUID), .BIT_WIDTH(64'd1)) And_39 (.in0(wire_48), .in1(wire_39), .out(wire_20));
  TC_Halt # (.UUID(64'd1474802306642119463 ^ UUID), .HALT_MESSAGE("End of file reached!")) Halt_40 (.clk(clk), .rst(rst), .en(wire_32));
  TC_Halt # (.UUID(64'd3727559317572521050 ^ UUID), .HALT_MESSAGE("Found crossing")) Halt_41 (.clk(clk), .rst(rst), .en(1'd0));
  TC_And3 # (.UUID(64'd3134744527415087055 ^ UUID), .BIT_WIDTH(64'd1)) And3_42 (.in0(wire_0), .in1(wire_20), .in2(wire_12), .out(wire_32));
  TC_FileLoader # (.UUID(64'd3429124062269983960 ^ UUID), .DEFAULT_FILE_NAME("day3_test_2")) FileLoader_43 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_25), .out(wire_5_1));
  TC_FileLoader # (.UUID(64'd1473616339079632962 ^ UUID), .DEFAULT_FILE_NAME("day3_test_3")) FileLoader_44 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_25), .out(wire_5_3));
  TC_Halt # (.UUID(64'd2886596719389344914 ^ UUID), .HALT_MESSAGE("Adder overflow! (PositionAdder)")) Halt_45 (.clk(clk), .rst(rst), .en(1'd0));
  TC_DelayLine # (.UUID(64'd4084865240337909835 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_46 (.clk(clk), .rst(rst), .in(wire_18), .out(wire_50));
  TC_Counter # (.UUID(64'd1078548748747073918 ^ UUID), .BIT_WIDTH(64'd32), .count(32'd1)) Counter32_47 (.clk(clk), .rst(rst), .save(wire_24), .in(wire_51), .out(wire_14));
  TC_Mux # (.UUID(64'd1505105403550165448 ^ UUID), .BIT_WIDTH(64'd16)) Mux16_48 (.sel(wire_8), .in0(wire_13[15:0]), .in1(wire_1[15:0]), .out(wire_67));
  TC_Mux # (.UUID(64'd3012025827690671150 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_49 (.sel(wire_54), .in0(wire_13), .in1({{48{1'b0}}, wire_67 }), .out(wire_49));
  TC_DelayLine # (.UUID(64'd4321725562030923891 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_50 (.clk(clk), .rst(rst), .in(wire_34), .out(wire_13));
  TC_Constant # (.UUID(64'd1801593110111524660 ^ UUID), .BIT_WIDTH(64'd64), .value(64'hFFFFFFFFFFFFFFFF)) Constant64_51 (.out(wire_27));
  TC_Switch # (.UUID(64'd2129707110641163321 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_52 (.en(wire_57), .in(wire_27), .out(wire_34_1));
  TC_Switch # (.UUID(64'd3550382538366520995 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_53 (.en(wire_9), .in(wire_49), .out(wire_34_0));
  TC_DelayLine # (.UUID(64'd1099126945014138228 ^ UUID), .BIT_WIDTH(64'd64)) DelayLine64_54 (.clk(clk), .rst(rst), .in(wire_22), .out(wire_3));
  TC_LessU # (.UUID(64'd331889225750388357 ^ UUID), .BIT_WIDTH(64'd64)) LessU64_55 (.in0({{32{1'b0}}, wire_1 }), .in1(wire_13), .out(wire_8));
  TC_FileLoader # (.UUID(64'd784893077974596701 ^ UUID), .DEFAULT_FILE_NAME("day3_test_4")) FileLoader_56 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_25), .out(wire_5_4));
  TC_FileLoader # (.UUID(64'd224237426130976828 ^ UUID), .DEFAULT_FILE_NAME("day3_test_5")) FileLoader_57 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_25), .out(wire_5_5));
  TC_FileLoader # (.UUID(64'd4283039450414421346 ^ UUID), .DEFAULT_FILE_NAME("day3_test_6")) FileLoader_58 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_25), .out(wire_5_6));
  TC_FileLoader # (.UUID(64'd1657938444342303651 ^ UUID), .DEFAULT_FILE_NAME("day3_test_7")) FileLoader_59 (.clk(clk), .rst(rst), .en(1'd0), .address(wire_25), .out(wire_5_7));
  TC_NoteSound # (.UUID(64'd428366861129437171 ^ UUID)) NoteSound_60 (.clk(clk), .rst(rst), .command({{7{1'b0}}, wire_32 }), .note(8'd0), .pitch(8'd0));
  TC_Equal # (.UUID(64'd2258306651148961062 ^ UUID), .BIT_WIDTH(64'd64)) Equal64_61 (.in0({{32{1'b0}}, wire_1 }), .in1(wire_46), .out(wire_68));
  TC_Constant # (.UUID(64'd4013474236969664718 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h114)) Constant64_62 (.out(wire_46));
  TC_Halt # (.UUID(64'd3904806610885250207 ^ UUID), .HALT_MESSAGE("Debug halt")) Halt_63 (.clk(clk), .rst(rst), .en(wire_68));
  InputMananger # (.UUID(64'd280349663464583758 ^ UUID)) InputMananger_64 (.clk(clk), .rst(rst), .Main_8b(wire_58), .Offset(wire_62), .Output(wire_31), .NewLine(wire_44));
  QuickSave # (.UUID(64'd3964331221245691836 ^ UUID)) QuickSave_65 (.clk(clk), .rst(rst), .Value(wire_5), .\Number_(stored) (wire_37), .\Saved?_1 (wire_0), .\Saved?_2 (wire_56));
  ManhattanDistance # (.UUID(64'd4534475870914388036 ^ UUID)) ManhattanDistance_66 (.clk(clk), .rst(rst), .X(wire_59), .Y(wire_7), .Output(wire_1));
  CellRotator # (.UUID(64'd2988738449177159528 ^ UUID)) CellRotator_67 (.clk(clk), .rst(rst), .Tick(wire_20), .Input(wire_61), .Pos_2(wire_11), .Pos_1(wire_30), .Written());
  QuickSave # (.UUID(64'd3551179199781681902 ^ UUID)) QuickSave_68 (.clk(clk), .rst(rst), .Value({{63{1'b0}}, wire_44 }), .\Number_(stored) (wire_43), .\Saved?_1 (wire_47), .\Saved?_2 ());
  OnOrOff # (.UUID(64'd2880407376120648954 ^ UUID)) OnOrOff_69 (.clk(clk), .rst(rst), .Input(wire_65), .Output(wire_24));
  QuickSave # (.UUID(64'd4013860832325939171 ^ UUID)) QuickSave_70 (.clk(clk), .rst(rst), .Value({{32{1'b0}}, wire_10 }), .\Number_(stored) (wire_42), .\Saved?_1 (wire_39), .\Saved?_2 ());
  OnOrOff # (.UUID(64'd685402883028759750 ^ UUID)) OnOrOff_71 (.clk(clk), .rst(rst), .Input(wire_26), .Output(wire_19_1));
  OnOrOff # (.UUID(64'd2586521289870388092 ^ UUID)) OnOrOff_72 (.clk(clk), .rst(rst), .Input(wire_20), .Output(wire_19_0));
  PositionAdder # (.UUID(64'd1952379698983790479 ^ UUID)) PositionAdder_73 (.clk(clk), .rst(rst), .Current_Position(wire_50), .Move({{32{1'b0}}, wire_31 }), .overflow(wire_66), .New_Position(wire_18));
  PositionAdder # (.UUID(64'd549660374295142354 ^ UUID)) PositionAdder_74 (.clk(clk), .rst(rst), .Current_Position(wire_11), .Move({{32{1'b0}}, wire_31 }), .overflow(), .New_Position(wire_61));
  LineCrosserz_3 # (.UUID(64'd235678000759494782 ^ UUID)) LineCrosserz_3_75 (.clk(clk), .rst(rst), .L2End(wire_11), .L2Start(wire_30), .L1End(wire_22), .L1Start(wire_3), .Output_1(wire_54), .Output_2(wire_17));
  _64bz_toz_32b # (.UUID(64'd4074607966076726035 ^ UUID)) _64bz_toz_32b_76 (.clk(clk), .rst(rst), .Input(wire_3), .Output_1(wire_33), .Output_2(wire_63));
  _64bz_toz_32b # (.UUID(64'd3297953936306396081 ^ UUID)) _64bz_toz_32b_77 (.clk(clk), .rst(rst), .Input(wire_22), .Output_1(wire_15), .Output_2(wire_4));
  _64bz_toz_32b # (.UUID(64'd2799350786039608227 ^ UUID)) _64bz_toz_32b_78 (.clk(clk), .rst(rst), .Input(wire_30), .Output_1(wire_2), .Output_2(wire_23));
  _64bz_toz_32b # (.UUID(64'd4547022319690718172 ^ UUID)) _64bz_toz_32b_79 (.clk(clk), .rst(rst), .Input(wire_11), .Output_1(wire_40), .Output_2(wire_29));
  _64bz_toz_32b # (.UUID(64'd36584691338760372 ^ UUID)) _64bz_toz_32b_80 (.clk(clk), .rst(rst), .Input(wire_17), .Output_1(wire_7), .Output_2(wire_59));
  _64bz_toz_32b # (.UUID(64'd1683694981542803589 ^ UUID)) _64bz_toz_32b_81 (.clk(clk), .rst(rst), .Input(wire_50), .Output_1(wire_28), .Output_2(wire_38));
  NumberDisplayz_zmz_1rzm10d # (.UUID(64'd1558355514723882557 ^ UUID)) NumberDisplayz_zmz_1rzm10d_82 (.clk(clk), .rst(rst), .Input(wire_38));
  NumberDisplayz_zmz_1rzm10d # (.UUID(64'd1342504794432391415 ^ UUID)) NumberDisplayz_zmz_1rzm10d_83 (.clk(clk), .rst(rst), .Input(wire_28));
  TC_Switch # (.UUID(64'd2241906331493591448 ^ UUID), .BIT_WIDTH(64'd64)) Switch64_84 (.en(wire_16), .in(wire_5), .out(wire_58));

  wire [0:0] wire_0;
  wire [31:0] wire_1;
  wire [31:0] wire_2;
  wire [63:0] wire_3;
  wire [31:0] wire_4;
  wire [63:0] wire_5;
  wire [63:0] wire_5_0;
  wire [63:0] wire_5_1;
  wire [63:0] wire_5_2;
  wire [63:0] wire_5_3;
  wire [63:0] wire_5_4;
  wire [63:0] wire_5_5;
  wire [63:0] wire_5_6;
  wire [63:0] wire_5_7;
  assign wire_5 = wire_5_0|wire_5_1|wire_5_2|wire_5_3|wire_5_4|wire_5_5|wire_5_6|wire_5_7;
  wire [0:0] wire_6;
  wire [31:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [31:0] wire_10;
  wire [63:0] wire_11;
  wire [0:0] wire_12;
  wire [63:0] wire_13;
  wire [31:0] wire_14;
  wire [31:0] wire_15;
  wire [0:0] wire_16;
  wire [63:0] wire_17;
  wire [63:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_19_0;
  wire [0:0] wire_19_1;
  assign wire_19 = wire_19_0|wire_19_1;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [63:0] wire_22;
  wire [31:0] wire_23;
  wire [0:0] wire_24;
  wire [63:0] wire_25;
  wire [0:0] wire_26;
  wire [63:0] wire_27;
  wire [31:0] wire_28;
  wire [31:0] wire_29;
  wire [63:0] wire_30;
  wire [31:0] wire_31;
  wire [0:0] wire_32;
  wire [31:0] wire_33;
  wire [63:0] wire_34;
  wire [63:0] wire_34_0;
  wire [63:0] wire_34_1;
  assign wire_34 = wire_34_0|wire_34_1;
  wire [63:0] wire_35;
  wire [0:0] wire_36;
  wire [63:0] wire_37;
  wire [31:0] wire_38;
  wire [0:0] wire_39;
  wire [31:0] wire_40;
  wire [63:0] wire_41;
  wire [63:0] wire_42;
  wire [63:0] wire_43;
  wire [0:0] wire_44;
  wire [63:0] wire_45;
  wire [63:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [63:0] wire_49;
  wire [63:0] wire_50;
  wire [31:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [63:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  wire [63:0] wire_58;
  wire [31:0] wire_59;
  wire [0:0] wire_60;
  wire [63:0] wire_61;
  wire [7:0] wire_62;
  wire [31:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [15:0] wire_67;
  wire [0:0] wire_68;

endmodule
